// ----------------------------------------------------------------------------
// LegUp High-Level Synthesis Tool Version 7.5 (http://legupcomputing.com)
// Copyright (c) 2015-2019 LegUp Computing Inc. All Rights Reserved.
// For technical issues, please contact: support@legupcomputing.com
// For general inquiries, please contact: info@legupcomputing.com
// Date: Fri Jun 26 12:00:36 2020
// ----------------------------------------------------------------------------
`define MEMORY_CONTROLLER_ADDR_SIZE 32
// This directory contains the memory initialization files generated by LegUp.
// This relative path is used by ModelSim and FPGA synthesis tool.
`define MEM_INIT_DIR "../mem_init/"

`timescale 1 ns / 1 ns
module top
(
	clk,
	reset,
	start,
	finish,
	return_val
);

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg  main_inst_clk;
reg  main_inst_reset;
reg  main_inst_start;
wire  main_inst_finish;
wire [31:0] main_inst_return_val;
reg  main_inst_finish_reg;
reg [31:0] main_inst_return_val_reg;


main main_inst (
	.clk (main_inst_clk),
	.reset (main_inst_reset),
	.start (main_inst_start),
	.finish (main_inst_finish),
	.return_val (main_inst_return_val)
);



always @(*) begin
	main_inst_clk = clk;
end
always @(*) begin
	main_inst_reset = reset;
end
always @(*) begin
	main_inst_start = start;
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_finish_reg <= 1'd0;
	end
	if (main_inst_finish) begin
		main_inst_finish_reg <= 1'd1;
	end
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_return_val_reg <= 0;
	end
	if (main_inst_finish) begin
		main_inst_return_val_reg <= main_inst_return_val;
	end
end
always @(*) begin
	finish = main_inst_finish;
end
always @(*) begin
	return_val = main_inst_return_val;
end

endmodule
`timescale 1 ns / 1 ns
module main
(
	clk,
	reset,
	start,
	finish,
	return_val
);

parameter [7:0] LEGUP_0 = 8'd0;
parameter [7:0] LEGUP_F_main_BB_while_body_lr_ph_1 = 8'd1;
parameter [7:0] LEGUP_F_main_BB_while_body_i_2 = 8'd2;
parameter [7:0] LEGUP_F_main_BB_while_body_i_3 = 8'd3;
parameter [7:0] LEGUP_F_main_BB_legup_memset_4_exit_4 = 8'd4;
parameter [7:0] LEGUP_F_main_BB_legup_memset_4_exit_5 = 8'd5;
parameter [7:0] LEGUP_F_main_BB_legup_memset_4_exit_6 = 8'd6;
parameter [7:0] LEGUP_F_main_BB_legup_memset_4_exit_7 = 8'd7;
parameter [7:0] LEGUP_F_main_BB_legup_memset_4_exit_8 = 8'd8;
parameter [7:0] LEGUP_F_main_BB_legup_memset_4_exit_9 = 8'd9;
parameter [7:0] LEGUP_F_main_BB_legup_memset_4_exit_10 = 8'd10;
parameter [7:0] LEGUP_F_main_BB_legup_memset_4_exit_11 = 8'd11;
parameter [7:0] LEGUP_F_main_BB_legup_memset_4_exit_12 = 8'd12;
parameter [7:0] LEGUP_F_main_BB_legup_memset_4_exit_13 = 8'd13;
parameter [7:0] LEGUP_F_main_BB_legup_memset_4_exit_14 = 8'd14;
parameter [7:0] LEGUP_F_main_BB_while_body_15 = 8'd15;
parameter [7:0] LEGUP_F_main_BB_while_body_16 = 8'd16;
parameter [7:0] LEGUP_F_main_BB_NodeBlock11_17 = 8'd17;
parameter [7:0] LEGUP_F_main_BB_NodeBlock9_18 = 8'd18;
parameter [7:0] LEGUP_F_main_BB_LeafBlock7_19 = 8'd19;
parameter [7:0] LEGUP_F_main_BB_LeafBlock5_20 = 8'd20;
parameter [7:0] LEGUP_F_main_BB_LeafBlock3_21 = 8'd21;
parameter [7:0] LEGUP_F_main_BB_NodeBlock_22 = 8'd22;
parameter [7:0] LEGUP_F_main_BB_LeafBlock1_23 = 8'd23;
parameter [7:0] LEGUP_F_main_BB_LeafBlock_24 = 8'd24;
parameter [7:0] LEGUP_F_main_BB_sw_bb_i_25 = 8'd25;
parameter [7:0] LEGUP_F_main_BB_if_then_i_26 = 8'd26;
parameter [7:0] LEGUP_F_main_BB_if_else_i_27 = 8'd27;
parameter [7:0] LEGUP_F_main_BB_sw_bb40_i_28 = 8'd28;
parameter [7:0] LEGUP_F_main_BB_if_then44_i_29 = 8'd29;
parameter [7:0] LEGUP_F_main_BB_if_else62_i_30 = 8'd30;
parameter [7:0] LEGUP_F_main_BB_sw_bb84_i_31 = 8'd31;
parameter [7:0] LEGUP_F_main_BB_if_then88_i_32 = 8'd32;
parameter [7:0] LEGUP_F_main_BB_sw_epilog_thread242_i_33 = 8'd33;
parameter [7:0] LEGUP_F_main_BB_sw_bb118_i_34 = 8'd34;
parameter [7:0] LEGUP_F_main_BB_sw_default_i_35 = 8'd35;
parameter [7:0] LEGUP_F_main_BB_if_then126_i_36 = 8'd36;
parameter [7:0] LEGUP_F_main_BB_if_else131_i_37 = 8'd37;
parameter [7:0] LEGUP_F_main_BB_NodeBlock24_38 = 8'd38;
parameter [7:0] LEGUP_F_main_BB_NodeBlock22_39 = 8'd39;
parameter [7:0] LEGUP_F_main_BB_LeafBlock20_40 = 8'd40;
parameter [7:0] LEGUP_F_main_BB_LeafBlock18_41 = 8'd41;
parameter [7:0] LEGUP_F_main_BB_LeafBlock16_42 = 8'd42;
parameter [7:0] LEGUP_F_main_BB_sw_default142_i_43 = 8'd43;
parameter [7:0] LEGUP_F_main_BB_NodeBlock43_44 = 8'd44;
parameter [7:0] LEGUP_F_main_BB_NodeBlock41_45 = 8'd45;
parameter [7:0] LEGUP_F_main_BB_NodeBlock39_46 = 8'd46;
parameter [7:0] LEGUP_F_main_BB_LeafBlock37_47 = 8'd47;
parameter [7:0] LEGUP_F_main_BB_LeafBlock35_48 = 8'd48;
parameter [7:0] LEGUP_F_main_BB_LeafBlock33_49 = 8'd49;
parameter [7:0] LEGUP_F_main_BB_NodeBlock31_50 = 8'd50;
parameter [7:0] LEGUP_F_main_BB_LeafBlock29_51 = 8'd51;
parameter [7:0] LEGUP_F_main_BB_LeafBlock27_52 = 8'd52;
parameter [7:0] LEGUP_F_main_BB_sw_default148_i_53 = 8'd53;
parameter [7:0] LEGUP_F_main_BB_NodeBlock78_54 = 8'd54;
parameter [7:0] LEGUP_F_main_BB_NodeBlock76_55 = 8'd55;
parameter [7:0] LEGUP_F_main_BB_NodeBlock74_56 = 8'd56;
parameter [7:0] LEGUP_F_main_BB_NodeBlock72_57 = 8'd57;
parameter [7:0] LEGUP_F_main_BB_LeafBlock70_58 = 8'd58;
parameter [7:0] LEGUP_F_main_BB_LeafBlock68_59 = 8'd59;
parameter [7:0] LEGUP_F_main_BB_LeafBlock66_60 = 8'd60;
parameter [7:0] LEGUP_F_main_BB_NodeBlock64_61 = 8'd61;
parameter [7:0] LEGUP_F_main_BB_LeafBlock62_62 = 8'd62;
parameter [7:0] LEGUP_F_main_BB_LeafBlock60_63 = 8'd63;
parameter [7:0] LEGUP_F_main_BB_NodeBlock58_64 = 8'd64;
parameter [7:0] LEGUP_F_main_BB_NodeBlock56_65 = 8'd65;
parameter [7:0] LEGUP_F_main_BB_LeafBlock54_66 = 8'd66;
parameter [7:0] LEGUP_F_main_BB_LeafBlock52_67 = 8'd67;
parameter [7:0] LEGUP_F_main_BB_NodeBlock50_68 = 8'd68;
parameter [7:0] LEGUP_F_main_BB_LeafBlock48_69 = 8'd69;
parameter [7:0] LEGUP_F_main_BB_LeafBlock46_70 = 8'd70;
parameter [7:0] LEGUP_F_main_BB_NodeBlock89_71 = 8'd71;
parameter [7:0] LEGUP_F_main_BB_NodeBlock87_72 = 8'd72;
parameter [7:0] LEGUP_F_main_BB_LeafBlock85_73 = 8'd73;
parameter [7:0] LEGUP_F_main_BB_LeafBlock83_74 = 8'd74;
parameter [7:0] LEGUP_F_main_BB_LeafBlock81_75 = 8'd75;
parameter [7:0] LEGUP_F_main_BB_NodeBlock96_76 = 8'd76;
parameter [7:0] LEGUP_F_main_BB_LeafBlock94_77 = 8'd77;
parameter [7:0] LEGUP_F_main_BB_LeafBlock92_78 = 8'd78;
parameter [7:0] LEGUP_F_main_BB_sw_default13_i_79 = 8'd79;
parameter [7:0] LEGUP_F_main_BB_sw_default16_i_80 = 8'd80;
parameter [7:0] LEGUP_F_main_BB_NodeBlock115_81 = 8'd81;
parameter [7:0] LEGUP_F_main_BB_NodeBlock113_82 = 8'd82;
parameter [7:0] LEGUP_F_main_BB_NodeBlock111_83 = 8'd83;
parameter [7:0] LEGUP_F_main_BB_LeafBlock109_84 = 8'd84;
parameter [7:0] LEGUP_F_main_BB_LeafBlock109_sw_default31_i_crit_edge_85 = 8'd85;
parameter [7:0] LEGUP_F_main_BB_NodeBlock107_86 = 8'd86;
parameter [7:0] LEGUP_F_main_BB_NodeBlock105_87 = 8'd87;
parameter [7:0] LEGUP_F_main_BB_NodeBlock103_88 = 8'd88;
parameter [7:0] LEGUP_F_main_BB_NodeBlock101_89 = 8'd89;
parameter [7:0] LEGUP_F_main_BB_LeafBlock99_90 = 8'd90;
parameter [7:0] LEGUP_F_main_BB_LeafBlock99_sw_default31_i_crit_edge_91 = 8'd91;
parameter [7:0] LEGUP_F_main_BB_NodeBlock122_92 = 8'd92;
parameter [7:0] LEGUP_F_main_BB_LeafBlock120_93 = 8'd93;
parameter [7:0] LEGUP_F_main_BB_LeafBlock118_94 = 8'd94;
parameter [7:0] LEGUP_F_main_BB_sw_default29_i_95 = 8'd95;
parameter [7:0] LEGUP_F_main_BB_sw_default31_i_96 = 8'd96;
parameter [7:0] LEGUP_F_main_BB_sw_default48_i_97 = 8'd97;
parameter [7:0] LEGUP_F_main_BB_switch_lookup_i_98 = 8'd98;
parameter [7:0] LEGUP_F_main_BB_switch_lookup_i_99 = 8'd99;
parameter [7:0] LEGUP_F_main_BB_switch_lookup54_i_100 = 8'd100;
parameter [7:0] LEGUP_F_main_BB_switch_lookup54_i_101 = 8'd101;
parameter [7:0] LEGUP_F_main_BB_aluDecode_exit_102 = 8'd102;
parameter [7:0] LEGUP_F_main_BB_aluDecode_exit_103 = 8'd103;
parameter [7:0] LEGUP_F_main_BB_if_else_104 = 8'd104;
parameter [7:0] LEGUP_F_main_BB_if_else_105 = 8'd105;
parameter [7:0] LEGUP_F_main_BB_NodeBlock175_106 = 8'd106;
parameter [7:0] LEGUP_F_main_BB_NodeBlock173_107 = 8'd107;
parameter [7:0] LEGUP_F_main_BB_NodeBlock171_108 = 8'd108;
parameter [7:0] LEGUP_F_main_BB_NodeBlock169_109 = 8'd109;
parameter [7:0] LEGUP_F_main_BB_NodeBlock167_110 = 8'd110;
parameter [7:0] LEGUP_F_main_BB_LeafBlock165_111 = 8'd111;
parameter [7:0] LEGUP_F_main_BB_NodeBlock163_112 = 8'd112;
parameter [7:0] LEGUP_F_main_BB_NodeBlock161_113 = 8'd113;
parameter [7:0] LEGUP_F_main_BB_LeafBlock159_114 = 8'd114;
parameter [7:0] LEGUP_F_main_BB_NodeBlock157_115 = 8'd115;
parameter [7:0] LEGUP_F_main_BB_NodeBlock155_116 = 8'd116;
parameter [7:0] LEGUP_F_main_BB_NodeBlock153_117 = 8'd117;
parameter [7:0] LEGUP_F_main_BB_NodeBlock151_118 = 8'd118;
parameter [7:0] LEGUP_F_main_BB_NodeBlock149_119 = 8'd119;
parameter [7:0] LEGUP_F_main_BB_NodeBlock147_120 = 8'd120;
parameter [7:0] LEGUP_F_main_BB_NodeBlock145_121 = 8'd121;
parameter [7:0] LEGUP_F_main_BB_NodeBlock143_122 = 8'd122;
parameter [7:0] LEGUP_F_main_BB_NodeBlock141_123 = 8'd123;
parameter [7:0] LEGUP_F_main_BB_NodeBlock139_124 = 8'd124;
parameter [7:0] LEGUP_F_main_BB_NodeBlock137_125 = 8'd125;
parameter [7:0] LEGUP_F_main_BB_NodeBlock135_126 = 8'd126;
parameter [7:0] LEGUP_F_main_BB_NodeBlock133_127 = 8'd127;
parameter [7:0] LEGUP_F_main_BB_NodeBlock131_128 = 8'd128;
parameter [7:0] LEGUP_F_main_BB_NodeBlock129_129 = 8'd129;
parameter [7:0] LEGUP_F_main_BB_NodeBlock127_130 = 8'd130;
parameter [7:0] LEGUP_F_main_BB_LeafBlock125_131 = 8'd131;
parameter [7:0] LEGUP_F_main_BB_sw_bb1_i_132 = 8'd132;
parameter [7:0] LEGUP_F_main_BB_sw_bb5_i_133 = 8'd133;
parameter [7:0] LEGUP_F_main_BB_sw_bb9_i_134 = 8'd134;
parameter [7:0] LEGUP_F_main_BB_sw_bb13_i_135 = 8'd135;
parameter [7:0] LEGUP_F_main_BB_sw_bb17_i_136 = 8'd136;
parameter [7:0] LEGUP_F_main_BB_sw_bb22_i_137 = 8'd137;
parameter [7:0] LEGUP_F_main_BB_sw_bb31_i_138 = 8'd138;
parameter [7:0] LEGUP_F_main_BB_sw_bb37_i_139 = 8'd139;
parameter [7:0] LEGUP_F_main_BB_sw_bb42_i_140 = 8'd140;
parameter [7:0] LEGUP_F_main_BB_sw_bb49_i_141 = 8'd141;
parameter [7:0] LEGUP_F_main_BB_sw_bb54_i_142 = 8'd142;
parameter [7:0] LEGUP_F_main_BB_sw_bb60_i_143 = 8'd143;
parameter [7:0] LEGUP_F_main_BB_sw_bb65_i_144 = 8'd144;
parameter [7:0] LEGUP_F_main_BB_sw_bb65_i_145 = 8'd145;
parameter [7:0] LEGUP_F_main_BB_sw_bb73_i_146 = 8'd146;
parameter [7:0] LEGUP_F_main_BB_sw_bb83_i_147 = 8'd147;
parameter [7:0] LEGUP_F_main_BB_sw_bb88_i_148 = 8'd148;
parameter [7:0] LEGUP_F_main_BB_sw_bb97_i_149 = 8'd149;
parameter [7:0] LEGUP_F_main_BB_sw_bb106_i_150 = 8'd150;
parameter [7:0] LEGUP_F_main_BB_sw_bb115_i_151 = 8'd151;
parameter [7:0] LEGUP_F_main_BB_sw_bb124_i_152 = 8'd152;
parameter [7:0] LEGUP_F_main_BB_sw_bb133_i_153 = 8'd153;
parameter [7:0] LEGUP_F_main_BB_alu_exit_154 = 8'd154;
parameter [7:0] LEGUP_F_main_BB_if_then38_155 = 8'd155;
parameter [7:0] LEGUP_F_main_BB_if_then38_156 = 8'd156;
parameter [7:0] LEGUP_F_main_BB_if_then38_157 = 8'd157;
parameter [7:0] LEGUP_F_main_BB_if_end42_158 = 8'd158;
parameter [7:0] LEGUP_F_main_BB_if_then47_159 = 8'd159;
parameter [7:0] LEGUP_F_main_BB_if_then47_160 = 8'd160;
parameter [7:0] LEGUP_F_main_BB_if_then47_161 = 8'd161;
parameter [7:0] LEGUP_F_main_BB_if_else51_162 = 8'd162;
parameter [7:0] LEGUP_F_main_BB_if_then56_163 = 8'd163;
parameter [7:0] LEGUP_F_main_BB_if_then56_164 = 8'd164;
parameter [7:0] LEGUP_F_main_BB_if_end61_165 = 8'd165;
parameter [7:0] LEGUP_F_main_BB_if_then_i1_166 = 8'd166;
parameter [7:0] LEGUP_F_main_BB_if_then8_i_167 = 8'd167;
parameter [7:0] LEGUP_F_main_BB_if_else_i2_168 = 8'd168;
parameter [7:0] LEGUP_F_main_BB_if_then13_i_169 = 8'd169;
parameter [7:0] LEGUP_F_main_BB_if_else15_i_170 = 8'd170;
parameter [7:0] LEGUP_F_main_BB_if_else18_i_171 = 8'd171;
parameter [7:0] LEGUP_F_main_BB_addressCalculator_exit_172 = 8'd172;
parameter [7:0] LEGUP_F_main_BB_if_end61_while_body_crit_edge_173 = 8'd173;
parameter [7:0] LEGUP_F_main_BB_if_end61_while_body_crit_edge_174 = 8'd174;
parameter [7:0] LEGUP_F_main_BB_while_end_175 = 8'd175;
parameter [7:0] LEGUP_F_main_BB_while_end_176 = 8'd176;

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg [7:0] cur_state/* synthesis syn_encoding="onehot" */;
reg [7:0] next_state;
wire  fsm_stall;
reg [5:0] main_while_body_i_indvar;
reg [5:0] main_while_body_i_indvar_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_while_body_i_s_010_i;
reg [6:0] main_while_body_i_0;
reg [6:0] main_while_body_i_0_reg;
reg  main_while_body_i_exitcond1;
reg  main_while_body_i_exitcond1_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx1;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx2;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx2_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx3;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx3_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx4;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx4_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx5;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx5_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx6;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx6_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx7;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx7_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx8;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx8_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx9;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx9_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx10;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx10_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx11;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx11_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx12;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx12_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx13;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx13_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx14;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx14_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx15;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx15_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx16;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx16_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx17;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx17_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx18;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx18_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx19;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx19_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx22;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_legup_memset_4_exit_arrayidx22_reg;
reg [31:0] main_while_body_1;
reg [31:0] main_while_body_1_reg;
reg [31:0] main_while_body_nextInst_099;
reg [31:0] main_while_body_nextInst_099_reg;
reg [4:0] main_while_body_bit_select44;
reg [4:0] main_while_body_bit_select42;
reg [2:0] main_while_body_bit_select39;
reg [6:0] main_while_body_bit_select37;
reg [9:0] main_while_body_bit_select32;
reg [9:0] main_while_body_bit_select32_reg;
reg [3:0] main_while_body_bit_select30;
reg [3:0] main_while_body_bit_select30_reg;
reg  main_while_body_bit_select29;
reg  main_while_body_bit_select29_reg;
reg [7:0] main_while_body_bit_select28;
reg [7:0] main_while_body_bit_select28_reg;
reg  main_while_body_bit_select25;
reg  main_while_body_bit_select25_reg;
reg [3:0] main_while_body_bit_select24;
reg [3:0] main_while_body_bit_select24_reg;
reg [4:0] main_while_body_bit_select23;
reg [4:0] main_while_body_bit_select23_reg;
reg [4:0] main_while_body_bit_select21;
reg [4:0] main_while_body_bit_select21_reg;
reg [5:0] main_while_body_bit_select20;
reg [5:0] main_while_body_bit_select20_reg;
reg [19:0] main_while_body_bit_select17;
reg [19:0] main_while_body_bit_select17_reg;
reg  main_while_body_bit_select16;
reg  main_while_body_bit_select16_reg;
reg [10:0] main_while_body_bit_select13;
reg [10:0] main_while_body_bit_select13_reg;
reg [31:0] main_while_body_bit_concat45;
reg [31:0] main_while_body_bit_concat45_reg;
reg [31:0] main_while_body_bit_concat43;
reg [31:0] main_while_body_bit_concat43_reg;
reg [31:0] main_while_body_bit_concat41;
reg [31:0] main_while_body_bit_concat41_reg;
reg [6:0] main_while_body_shr6_i;
reg [6:0] main_while_body_shr6_i_reg;
reg [31:0] main_while_body_bit_concat40;
reg [31:0] main_while_body_bit_concat40_reg;
reg [31:0] main_while_body_bit_concat38;
reg [31:0] main_while_body_bit_concat38_reg;
reg  main_while_body_Pivot14;
reg  main_while_body_Pivot14_reg;
reg  main_NodeBlock11_Pivot12;
reg  main_NodeBlock9_Pivot10;
reg  main_LeafBlock7_SwitchLeaf8;
reg  main_LeafBlock5_SwitchLeaf6;
reg  main_LeafBlock3_SwitchLeaf4;
reg  main_NodeBlock_Pivot;
reg  main_LeafBlock1_SwitchLeaf2;
reg  main_LeafBlock_SwitchLeaf;
reg [1:0] main_sw_bb_i_shr13_i;
reg  main_sw_bb_i_bit_select34;
reg  main_sw_bb_i_bit_select34_reg;
reg  main_sw_bb_i_cmp_i;
reg [31:0] main_if_then_i_bit_concat36;
reg [31:0] main_if_else_i_bit_concat35;
reg [1:0] main_sw_bb40_i_shr42_i;
reg  main_sw_bb40_i_bit_select27;
reg  main_sw_bb40_i_bit_select27_reg;
reg  main_sw_bb40_i_cmp43_i;
reg [31:0] main_if_then44_i_bit_concat33;
reg [31:0] main_if_else62_i_bit_concat31;
reg [1:0] main_sw_bb84_i_shr86_i;
reg  main_sw_bb84_i_bit_select19;
reg  main_sw_bb84_i_bit_select19_reg;
reg  main_sw_bb84_i_cmp87_i;
reg [31:0] main_if_then88_i_bit_concat26;
reg [31:0] main_sw_epilog_thread242_i_bit_concat22;
reg [31:0] main_sw_bb118_i_bit_concat18;
reg [31:0] main_if_then126_i_bit_concat15;
reg [31:0] main_if_else131_i_bit_concat14;
reg [31:0] main_NodeBlock24_results_sroa_14_0_i;
reg [31:0] main_NodeBlock24_results_sroa_14_0_i_reg;
reg  main_NodeBlock24_Pivot25;
reg  main_NodeBlock22_Pivot23;
reg  main_LeafBlock20_SwitchLeaf21;
reg  main_LeafBlock18_SwitchLeaf19;
reg  main_LeafBlock16_SwitchLeaf17;
reg [31:0] main_sw_default142_i_results_sroa_14_0243_i;
reg [31:0] main_sw_default142_i_results_sroa_14_0243_i_reg;
reg [31:0] main_NodeBlock43_results_sroa_14_0241_i;
reg [31:0] main_NodeBlock43_results_sroa_14_0241_i_reg;
reg  main_NodeBlock43_results_sroa_23_0_i;
reg  main_NodeBlock43_results_sroa_23_0_i_reg;
reg  main_NodeBlock43_Pivot44;
reg  main_NodeBlock41_Pivot42;
reg  main_LeafBlock37_SwitchLeaf38;
reg  main_LeafBlock35_SwitchLeaf36;
reg  main_LeafBlock33_SwitchLeaf34;
reg  main_NodeBlock31_Pivot32;
reg  main_LeafBlock29_SwitchLeaf30;
reg  main_LeafBlock27_SwitchLeaf28;
reg [16:0] main_sw_default148_i_results_sroa_28_0249_i;
reg [16:0] main_sw_default148_i_results_sroa_28_0249_i_reg;
reg  main_sw_default148_i_results_sroa_23_0247_i;
reg  main_sw_default148_i_results_sroa_23_0247_i_reg;
reg [31:0] main_sw_default148_i_results_sroa_14_0241245_i;
reg [31:0] main_sw_default148_i_results_sroa_14_0241245_i_reg;
reg [16:0] main_NodeBlock78_results_sroa_28_0248_i;
reg [16:0] main_NodeBlock78_results_sroa_28_0248_i_reg;
reg  main_NodeBlock78_results_sroa_23_0246_i;
reg  main_NodeBlock78_results_sroa_23_0246_i_reg;
reg [31:0] main_NodeBlock78_results_sroa_14_0241244_i;
reg [31:0] main_NodeBlock78_results_sroa_14_0241244_i_reg;
reg [8:0] main_NodeBlock78_results_sroa_26_0_i;
reg [8:0] main_NodeBlock78_results_sroa_26_0_i_reg;
reg  main_NodeBlock78_bit_select3;
reg  main_NodeBlock78_bit_select3_reg;
reg  main_NodeBlock78_bit_select1;
reg  main_NodeBlock78_bit_select1_reg;
reg  main_NodeBlock78_Pivot79;
reg  main_NodeBlock76_Pivot77;
reg  main_NodeBlock74_Pivot75;
reg  main_NodeBlock72_Pivot73;
reg  main_LeafBlock70_SwitchLeaf71;
reg  main_LeafBlock68_SwitchLeaf69;
reg  main_LeafBlock66_SwitchLeaf67;
reg  main_LeafBlock62_SwitchLeaf63;
reg  main_LeafBlock60_SwitchLeaf61;
reg  main_NodeBlock58_Pivot59;
reg  main_NodeBlock56_Pivot57;
reg  main_LeafBlock54_SwitchLeaf55;
reg  main_LeafBlock52_SwitchLeaf53;
reg  main_NodeBlock50_Pivot51;
reg  main_LeafBlock48_SwitchLeaf49;
reg  main_LeafBlock46_SwitchLeaf47;
reg  main_NodeBlock89_Pivot90;
reg  main_NodeBlock87_Pivot88;
reg  main_LeafBlock85_SwitchLeaf86;
reg  main_LeafBlock83_SwitchLeaf84;
reg  main_LeafBlock81_SwitchLeaf82;
reg  main_NodeBlock96_Pivot97;
reg  main_LeafBlock94_SwitchLeaf95;
reg  main_LeafBlock92_SwitchLeaf93;
reg  main_NodeBlock115_Pivot116;
reg  main_NodeBlock113_Pivot114;
reg  main_NodeBlock111_Pivot112;
reg  main_NodeBlock107_Pivot108;
reg  main_NodeBlock105_Pivot106;
reg  main_NodeBlock103_Pivot104;
reg [2:0] main_NodeBlock103_1;
reg  main_NodeBlock101_Pivot102;
reg  main_NodeBlock122_Pivot123;
reg  main_LeafBlock120_SwitchLeaf121;
reg  main_LeafBlock118_SwitchLeaf119;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_switch_lookup_i_switch_gep_i;
reg [31:0] main_switch_lookup_i_switch_load_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_switch_lookup54_i_switch_gep56_i;
reg [31:0] main_switch_lookup54_i_switch_load57_i;
reg [15:0] main_aluDecode_exit_results_sroa_37_0_i6;
reg [15:0] main_aluDecode_exit_results_sroa_37_0_i6_reg;
reg [31:0] main_aluDecode_exit_results_sroa_31_0250_i4;
reg [31:0] main_aluDecode_exit_results_sroa_31_0250_i4_reg;
reg [15:0] main_aluDecode_exit_results_sroa_34_0252_i2;
reg [15:0] main_aluDecode_exit_results_sroa_34_0252_i2_reg;
reg [31:0] main_aluDecode_exit_call13;
reg [31:0] main_aluDecode_exit_call13_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_aluDecode_exit_arrayidx24;
reg [31:0] main_aluDecode_exit_2;
reg [31:0] main_aluDecode_exit_2_reg;
reg  main_aluDecode_exit_tobool;
reg  main_aluDecode_exit_tobool_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_else_arrayidx27;
reg [31:0] main_if_else_3;
reg [31:0] main_NodeBlock175_aluB_0;
reg [31:0] main_NodeBlock175_aluB_0_reg;
reg  main_NodeBlock175_Pivot176;
reg  main_NodeBlock173_Pivot174;
reg  main_NodeBlock171_Pivot172;
reg  main_NodeBlock169_Pivot170;
reg  main_NodeBlock167_Pivot168;
reg  main_LeafBlock165_SwitchLeaf166;
reg  main_NodeBlock163_Pivot164;
reg  main_NodeBlock161_Pivot162;
reg  main_LeafBlock159_SwitchLeaf160;
reg  main_NodeBlock157_Pivot158;
reg  main_NodeBlock155_Pivot156;
reg  main_NodeBlock153_Pivot154;
reg  main_NodeBlock151_Pivot152;
reg  main_NodeBlock149_Pivot150;
reg  main_NodeBlock147_Pivot148;
reg  main_NodeBlock145_Pivot146;
reg  main_NodeBlock143_Pivot144;
reg  main_NodeBlock141_Pivot142;
reg  main_NodeBlock139_Pivot140;
reg  main_NodeBlock137_Pivot138;
reg  main_NodeBlock135_Pivot136;
reg  main_NodeBlock133_Pivot134;
reg  main_NodeBlock131_Pivot132;
reg  main_NodeBlock129_Pivot130;
reg  main_NodeBlock127_Pivot128;
reg  main_LeafBlock125_SwitchLeaf126;
reg [31:0] main_LeafBlock125_add_i4;
reg [31:0] main_LeafBlock125_add_i4_1;
reg [31:0] main_sw_bb1_i_sub_i;
reg [31:0] main_sw_bb5_i_and_i6;
reg [31:0] main_sw_bb9_i_or_i;
reg [31:0] main_sw_bb13_i_xor_i;
reg  main_sw_bb17_i_cmp_i7;
reg [31:0] main_sw_bb17_i_bit_concat12;
reg  main_sw_bb22_i_cmp23_i;
reg [31:0] main_sw_bb22_i_bit_concat11;
reg [31:0] main_sw_bb31_i_shr33_i;
reg [31:0] main_sw_bb37_i_shr38_i;
reg [31:0] main_sw_bb42_i_shr45_i;
reg [31:0] main_sw_bb49_i_shr50_i;
reg [31:0] main_sw_bb54_i_shl_i;
reg [31:0] main_sw_bb60_i_shl61_i;
reg [31:0] main_sw_bb65_i_mul_i;
reg [31:0] main_sw_bb73_i_add74_i;
reg [31:0] main_sw_bb83_i_add84_i;
reg  main_sw_bb88_i_cmp90_i;
reg [7:0] main_sw_bb88_i_bit_concat10;
reg  main_sw_bb97_i_not_cmp99_i;
reg [7:0] main_sw_bb97_i_bit_concat9;
reg  main_sw_bb106_i_cmp108_i;
reg [7:0] main_sw_bb106_i_bit_concat8;
reg  main_sw_bb115_i_not_cmp117_i;
reg [7:0] main_sw_bb115_i_bit_concat7;
reg  main_sw_bb124_i_cmp126_i;
reg [7:0] main_sw_bb124_i_bit_concat6;
reg  main_sw_bb133_i_not_cmp135_i;
reg [7:0] main_sw_bb133_i_bit_concat5;
reg [31:0] main_alu_exit_add79_i;
reg [31:0] main_alu_exit_add79_i_reg;
reg  main_alu_exit_tobool34;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then38_arrayidx40;
reg [31:0] main_if_then38_4;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then38_arrayidx41;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then38_arrayidx41_reg;
reg [31:0] main_if_end42_results_sroa_0_2_i16;
reg [31:0] main_if_end42_results_sroa_0_2_i16_reg;
reg [7:0] main_if_end42_results_sroa_53_6_i15;
reg [7:0] main_if_end42_results_sroa_53_6_i15_reg;
reg  main_if_end42_tobool43;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then47_arrayidx49;
reg [31:0] main_if_then47_5;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then47_arrayidx50;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then47_arrayidx50_reg;
reg  main_if_else51_tobool52;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then56_arrayidx59;
reg  main_if_end61_tobool63;
reg [31:0] main_if_end61_bit_concat4;
reg  main_if_end61_tobool66;
reg  main_if_end61_tobool66_reg;
reg [7:0] main_if_then_i1_bit_concat2;
reg  main_if_then_i1_tobool65;
reg [31:0] main_if_then8_i_add_i;
reg [31:0] main_if_then13_i_add14_i;
reg [30:0] main_if_then13_i_bit_select;
reg [31:0] main_if_then13_i_bit_concat;
reg [31:0] main_if_else15_i_add16_i;
reg [31:0] main_if_else18_i_add19_i;
reg [31:0] main_addressCalculator_exit_newPc_0_i;
reg [31:0] main_addressCalculator_exit_newPc_0_i_reg;
reg  main_addressCalculator_exit_cmp;
reg  main_addressCalculator_exit_cmp21;
reg  main_addressCalculator_exit_or_cond;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end61_while_body_crit_edge_arrayidx23_phi_;
reg [31:0] main_if_end61_while_body_crit_edge_pre100;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_while_end_arrayidx68_phi_trans_insert;
reg [31:0] main_while_end_pre;
reg [2:0] switch_table_address_a;
wire [31:0] switch_table_out_a;
wire [2:0] switch_table_address_b;
wire [31:0] switch_table_out_b;
reg [2:0] switch_table1_address_a;
wire [31:0] switch_table1_out_a;
wire [2:0] switch_table1_address_b;
wire [31:0] switch_table1_out_b;
reg [4:0] main_while_body_lr_ph_registers_address_a;
reg  main_while_body_lr_ph_registers_write_enable_a;
reg [31:0] main_while_body_lr_ph_registers_in_a;
wire [31:0] main_while_body_lr_ph_registers_out_a;
reg [9:0] main_while_body_lr_ph_instMemory_address_a;
reg  main_while_body_lr_ph_instMemory_write_enable_a;
reg [31:0] main_while_body_lr_ph_instMemory_in_a;
wire [31:0] main_while_body_lr_ph_instMemory_out_a;
reg [9:0] main_while_body_lr_ph_instMemory_address_b;
reg  main_while_body_lr_ph_instMemory_write_enable_b;
reg [31:0] main_while_body_lr_ph_instMemory_in_b;
wire [31:0] main_while_body_lr_ph_instMemory_out_b;
reg [12:0] main_while_body_lr_ph_memory_address_a;
reg  main_while_body_lr_ph_memory_write_enable_a;
reg [31:0] main_while_body_lr_ph_memory_in_a;
wire [31:0] main_while_body_lr_ph_memory_out_a;
wire [26:0] main_while_body_bit_concat45_bit_select_operand_0;
wire [26:0] main_while_body_bit_concat43_bit_select_operand_0;
wire [26:0] main_while_body_bit_concat41_bit_select_operand_0;
wire [28:0] main_while_body_bit_concat40_bit_select_operand_0;
wire [24:0] main_while_body_bit_concat38_bit_select_operand_0;
wire [20:0] main_if_then_i_bit_concat36_bit_select_operand_0;
wire  main_if_then_i_bit_concat36_bit_select_operand_6;
wire [17:0] main_if_else_i_bit_concat35_bit_select_operand_2;
wire  main_if_else_i_bit_concat35_bit_select_operand_6;
wire  main_if_else_i_bit_concat35_bit_select_operand_12;
wire [11:0] main_if_then44_i_bit_concat33_bit_select_operand_0;
wire  main_if_then44_i_bit_concat33_bit_select_operand_8;
wire [10:0] main_if_else62_i_bit_concat31_bit_select_operand_2;
wire  main_if_else62_i_bit_concat31_bit_select_operand_12;
wire [20:0] main_if_then88_i_bit_concat26_bit_select_operand_0;
wire  main_if_then88_i_bit_concat26_bit_select_operand_4;
wire [18:0] main_sw_epilog_thread242_i_bit_concat22_bit_select_operand_2;
wire  main_sw_epilog_thread242_i_bit_concat22_bit_select_operand_6;
wire [11:0] main_sw_bb118_i_bit_concat18_bit_select_operand_2;
wire [20:0] main_if_then126_i_bit_concat15_bit_select_operand_0;
wire [20:0] main_if_else131_i_bit_concat14_bit_select_operand_0;
wire [2:0] main_NodeBlock89_Pivot90_op1_temp;
wire [7:0] main_NodeBlock87_Pivot88_op1_temp;
wire [7:0] main_NodeBlock122_Pivot123_op1_temp;
wire [5:0] main_NodeBlock175_Pivot176_op1_temp;
wire [6:0] main_NodeBlock173_Pivot174_op1_temp;
wire [6:0] main_NodeBlock171_Pivot172_op1_temp;
wire [6:0] main_NodeBlock169_Pivot170_op1_temp;
wire [6:0] main_NodeBlock167_Pivot168_op1_temp;
wire [6:0] main_NodeBlock163_Pivot164_op1_temp;
wire [6:0] main_NodeBlock161_Pivot162_op1_temp;
wire [5:0] main_NodeBlock157_Pivot158_op1_temp;
wire [6:0] main_NodeBlock155_Pivot156_op1_temp;
wire [6:0] main_NodeBlock153_Pivot154_op1_temp;
wire [5:0] main_NodeBlock151_Pivot152_op1_temp;
wire [5:0] main_NodeBlock149_Pivot150_op1_temp;
wire [4:0] main_NodeBlock147_Pivot148_op1_temp;
wire [5:0] main_NodeBlock145_Pivot146_op1_temp;
wire [5:0] main_NodeBlock143_Pivot144_op1_temp;
wire [5:0] main_NodeBlock141_Pivot142_op1_temp;
wire [4:0] main_NodeBlock139_Pivot140_op1_temp;
wire [5:0] main_NodeBlock137_Pivot138_op1_temp;
wire [3:0] main_NodeBlock135_Pivot136_op1_temp;
wire [4:0] main_NodeBlock133_Pivot134_op1_temp;
wire [4:0] main_NodeBlock131_Pivot132_op1_temp;
wire [2:0] main_NodeBlock129_Pivot130_op1_temp;
wire [3:0] main_NodeBlock127_Pivot128_op1_temp;
wire [30:0] main_sw_bb17_i_bit_concat12_bit_select_operand_0;
wire [30:0] main_sw_bb22_i_bit_concat11_bit_select_operand_0;
reg  legup_mult_main_sw_bb65_i_mul_i_en;
reg [31:0] main_sw_bb65_i_mul_i_stage0_reg;
wire [6:0] main_sw_bb88_i_bit_concat10_bit_select_operand_0;
wire [6:0] main_sw_bb97_i_bit_concat9_bit_select_operand_0;
wire [6:0] main_sw_bb106_i_bit_concat8_bit_select_operand_0;
wire [6:0] main_sw_bb115_i_bit_concat7_bit_select_operand_0;
wire [6:0] main_sw_bb124_i_bit_concat6_bit_select_operand_0;
wire [6:0] main_sw_bb133_i_bit_concat5_bit_select_operand_0;
wire [14:0] main_if_end61_bit_concat4_bit_select_operand_0;
wire [15:0] main_if_end61_bit_concat4_bit_select_operand_4;
wire [6:0] main_if_then_i1_bit_concat2_bit_select_operand_0;
wire  main_if_then13_i_bit_concat_bit_select_operand_2;
wire [12:0] main_addressCalculator_exit_cmp21_op1_temp;



// @switch.table = private unnamed_addr constant [8 x i32] [i32 0, i32 11, i32 5, i32 6, i32 4, i32 9, i32 3, i32 2]
rom_dual_port switch_table (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( switch_table_address_a ),
	.q_a( switch_table_out_a ),
	.address_b( switch_table_address_b ),
	.q_b( switch_table_out_b )
);
defparam switch_table.width_a = 32;
defparam switch_table.widthad_a = 3;
defparam switch_table.numwords_a = 8;
defparam switch_table.width_b = 32;
defparam switch_table.widthad_b = 3;
defparam switch_table.numwords_b = 8;
defparam switch_table.latency = 1;
defparam switch_table.init_file = {`MEM_INIT_DIR, "switch_table.mif"};


// @switch.table1 = private unnamed_addr constant [8 x i32] [i32 20, i32 21, i32 31, i32 31, i32 23, i32 24, i32 25, i32 26]
rom_dual_port switch_table1 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( switch_table1_address_a ),
	.q_a( switch_table1_out_a ),
	.address_b( switch_table1_address_b ),
	.q_b( switch_table1_out_b )
);
defparam switch_table1.width_a = 32;
defparam switch_table1.widthad_a = 3;
defparam switch_table1.numwords_a = 8;
defparam switch_table1.width_b = 32;
defparam switch_table1.widthad_b = 3;
defparam switch_table1.numwords_b = 8;
defparam switch_table1.latency = 1;
defparam switch_table1.init_file = {`MEM_INIT_DIR, "switch_table1.mif"};


//   %registers = alloca [32 x i32], align 4, !MSB !96, !LSB !97, !extendFrom !96
ram_single_port_intel main_while_body_lr_ph_registers (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_while_body_lr_ph_registers_address_a ),
	.wren_a( main_while_body_lr_ph_registers_write_enable_a ),
	.data_a( main_while_body_lr_ph_registers_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_while_body_lr_ph_registers_out_a )
);
defparam main_while_body_lr_ph_registers.width_a = 32;
defparam main_while_body_lr_ph_registers.widthad_a = 5;
defparam main_while_body_lr_ph_registers.width_be_a = 4;
defparam main_while_body_lr_ph_registers.numwords_a = 32;
defparam main_while_body_lr_ph_registers.latency = 1;


//   %instMemory = alloca [1024 x i32], align 4, !MSB !96, !LSB !97, !extendFrom !96
ram_dual_port main_while_body_lr_ph_instMemory (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_while_body_lr_ph_instMemory_address_a ),
	.wren_a( main_while_body_lr_ph_instMemory_write_enable_a ),
	.data_a( main_while_body_lr_ph_instMemory_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_while_body_lr_ph_instMemory_out_a ),
	.address_b( main_while_body_lr_ph_instMemory_address_b ),
	.wren_b( main_while_body_lr_ph_instMemory_write_enable_b ),
	.data_b( main_while_body_lr_ph_instMemory_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_while_body_lr_ph_instMemory_out_b )
);
defparam main_while_body_lr_ph_instMemory.width_a = 32;
defparam main_while_body_lr_ph_instMemory.widthad_a = 10;
defparam main_while_body_lr_ph_instMemory.width_be_a = 4;
defparam main_while_body_lr_ph_instMemory.numwords_a = 1024;
defparam main_while_body_lr_ph_instMemory.width_b = 32;
defparam main_while_body_lr_ph_instMemory.widthad_b = 10;
defparam main_while_body_lr_ph_instMemory.width_be_b = 4;
defparam main_while_body_lr_ph_instMemory.numwords_b = 1024;
defparam main_while_body_lr_ph_instMemory.latency = 1;


//   %memory = alloca [8192 x i32], align 4, !MSB !96, !LSB !97, !extendFrom !96
ram_single_port_intel main_while_body_lr_ph_memory (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_while_body_lr_ph_memory_address_a ),
	.wren_a( main_while_body_lr_ph_memory_write_enable_a ),
	.data_a( main_while_body_lr_ph_memory_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_while_body_lr_ph_memory_out_a )
);
defparam main_while_body_lr_ph_memory.width_a = 32;
defparam main_while_body_lr_ph_memory.widthad_a = 13;
defparam main_while_body_lr_ph_memory.width_be_a = 4;
defparam main_while_body_lr_ph_memory.numwords_a = 8192;
defparam main_while_body_lr_ph_memory.latency = 1;

/* Unsynthesizable Statements */
/* synthesis translate_off */
always @(posedge clk)
	if (!fsm_stall) begin
	if ((cur_state == LEGUP_F_main_BB_while_end_176)) begin
		$write("%d\n", $signed(main_while_end_pre));
		// to fix quartus warning
		if (reset == 1'b0 && ^(main_while_end_pre) === 1'bX) finish <= 0;
	end
end
/* synthesis translate_on */
always @(posedge clk) begin
if (reset == 1'b1)
	cur_state <= LEGUP_0;
else if (!fsm_stall)
	cur_state <= next_state;
end

always @(*)
begin
next_state = cur_state;
case(cur_state)  /* synthesis parallel_case */
LEGUP_0:
	if ((fsm_stall == 1'd0) && (start == 1'd1))
		next_state = LEGUP_F_main_BB_while_body_lr_ph_1;
LEGUP_F_main_BB_LeafBlock109_84:
	if ((fsm_stall == 1'd0) && (1'd1 == 1'd1))
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
	else if ((fsm_stall == 1'd0) && (1'd1 == 1'd0))
		next_state = LEGUP_F_main_BB_LeafBlock109_sw_default31_i_crit_edge_85;
LEGUP_F_main_BB_LeafBlock109_sw_default31_i_crit_edge_85:
		next_state = LEGUP_F_main_BB_sw_default31_i_96;
LEGUP_F_main_BB_LeafBlock118_94:
	if ((fsm_stall == 1'd0) && (main_LeafBlock118_SwitchLeaf119 == 1'd1))
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock118_SwitchLeaf119 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default29_i_95;
LEGUP_F_main_BB_LeafBlock120_93:
	if ((fsm_stall == 1'd0) && (main_LeafBlock120_SwitchLeaf121 == 1'd1))
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock120_SwitchLeaf121 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default29_i_95;
LEGUP_F_main_BB_LeafBlock125_131:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_LeafBlock159_114:
	if ((fsm_stall == 1'd0) && (main_LeafBlock159_SwitchLeaf160 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb97_i_149;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock159_SwitchLeaf160 == 1'd0))
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_LeafBlock165_111:
	if ((fsm_stall == 1'd0) && (main_LeafBlock165_SwitchLeaf166 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb133_i_153;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock165_SwitchLeaf166 == 1'd0))
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_LeafBlock16_42:
	if ((fsm_stall == 1'd0) && (main_LeafBlock16_SwitchLeaf17 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock43_44;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock16_SwitchLeaf17 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default142_i_43;
LEGUP_F_main_BB_LeafBlock18_41:
	if ((fsm_stall == 1'd0) && (main_LeafBlock18_SwitchLeaf19 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_default148_i_53;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock18_SwitchLeaf19 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default142_i_43;
LEGUP_F_main_BB_LeafBlock1_23:
	if ((fsm_stall == 1'd0) && (main_LeafBlock1_SwitchLeaf2 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb84_i_31;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock1_SwitchLeaf2 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default_i_35;
LEGUP_F_main_BB_LeafBlock20_40:
	if ((fsm_stall == 1'd0) && (main_LeafBlock20_SwitchLeaf21 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock43_44;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock20_SwitchLeaf21 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default142_i_43;
LEGUP_F_main_BB_LeafBlock27_52:
	if ((fsm_stall == 1'd0) && (main_LeafBlock27_SwitchLeaf28 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock78_54;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock27_SwitchLeaf28 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default148_i_53;
LEGUP_F_main_BB_LeafBlock29_51:
	if ((fsm_stall == 1'd0) && (main_LeafBlock29_SwitchLeaf30 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock78_54;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock29_SwitchLeaf30 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default148_i_53;
LEGUP_F_main_BB_LeafBlock33_49:
	if ((fsm_stall == 1'd0) && (main_LeafBlock33_SwitchLeaf34 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock78_54;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock33_SwitchLeaf34 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default148_i_53;
LEGUP_F_main_BB_LeafBlock35_48:
	if ((fsm_stall == 1'd0) && (main_LeafBlock35_SwitchLeaf36 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock78_54;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock35_SwitchLeaf36 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default148_i_53;
LEGUP_F_main_BB_LeafBlock37_47:
	if ((fsm_stall == 1'd0) && (main_LeafBlock37_SwitchLeaf38 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock78_54;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock37_SwitchLeaf38 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default148_i_53;
LEGUP_F_main_BB_LeafBlock3_21:
	if ((fsm_stall == 1'd0) && (main_LeafBlock3_SwitchLeaf4 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb118_i_34;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock3_SwitchLeaf4 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default_i_35;
LEGUP_F_main_BB_LeafBlock46_70:
	if ((fsm_stall == 1'd0) && (main_LeafBlock46_SwitchLeaf47 == 1'd1))
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock46_SwitchLeaf47 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default48_i_97;
LEGUP_F_main_BB_LeafBlock48_69:
	if ((fsm_stall == 1'd0) && (main_LeafBlock48_SwitchLeaf49 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock115_81;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock48_SwitchLeaf49 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default48_i_97;
LEGUP_F_main_BB_LeafBlock52_67:
	if ((fsm_stall == 1'd0) && (main_LeafBlock52_SwitchLeaf53 == 1'd1))
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock52_SwitchLeaf53 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default48_i_97;
LEGUP_F_main_BB_LeafBlock54_66:
	if ((fsm_stall == 1'd0) && (main_LeafBlock54_SwitchLeaf55 == 1'd1))
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock54_SwitchLeaf55 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default48_i_97;
LEGUP_F_main_BB_LeafBlock5_20:
	if ((fsm_stall == 1'd0) && (main_LeafBlock5_SwitchLeaf6 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb_i_25;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock5_SwitchLeaf6 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default_i_35;
LEGUP_F_main_BB_LeafBlock60_63:
	if ((fsm_stall == 1'd0) && (main_LeafBlock60_SwitchLeaf61 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock89_71;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock60_SwitchLeaf61 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default48_i_97;
LEGUP_F_main_BB_LeafBlock62_62:
	if ((fsm_stall == 1'd0) && (main_LeafBlock62_SwitchLeaf63 == 1'd1))
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock62_SwitchLeaf63 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default48_i_97;
LEGUP_F_main_BB_LeafBlock66_60:
	if ((fsm_stall == 1'd0) && (main_LeafBlock66_SwitchLeaf67 == 1'd1))
		next_state = LEGUP_F_main_BB_switch_lookup54_i_100;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock66_SwitchLeaf67 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default48_i_97;
LEGUP_F_main_BB_LeafBlock68_59:
	if ((fsm_stall == 1'd0) && (main_LeafBlock68_SwitchLeaf69 == 1'd1))
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock68_SwitchLeaf69 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default48_i_97;
LEGUP_F_main_BB_LeafBlock70_58:
	if ((fsm_stall == 1'd0) && (main_LeafBlock70_SwitchLeaf71 == 1'd1))
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock70_SwitchLeaf71 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default48_i_97;
LEGUP_F_main_BB_LeafBlock7_19:
	if ((fsm_stall == 1'd0) && (main_LeafBlock7_SwitchLeaf8 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb40_i_28;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock7_SwitchLeaf8 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default_i_35;
LEGUP_F_main_BB_LeafBlock81_75:
	if ((fsm_stall == 1'd0) && (main_LeafBlock81_SwitchLeaf82 == 1'd1))
		next_state = LEGUP_F_main_BB_switch_lookup_i_98;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock81_SwitchLeaf82 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default16_i_80;
LEGUP_F_main_BB_LeafBlock83_74:
	if ((fsm_stall == 1'd0) && (main_LeafBlock83_SwitchLeaf84 == 1'd1))
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock83_SwitchLeaf84 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default16_i_80;
LEGUP_F_main_BB_LeafBlock85_73:
	if ((fsm_stall == 1'd0) && (main_LeafBlock85_SwitchLeaf86 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock96_76;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock85_SwitchLeaf86 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default16_i_80;
LEGUP_F_main_BB_LeafBlock92_78:
	if ((fsm_stall == 1'd0) && (main_LeafBlock92_SwitchLeaf93 == 1'd1))
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock92_SwitchLeaf93 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default13_i_79;
LEGUP_F_main_BB_LeafBlock94_77:
	if ((fsm_stall == 1'd0) && (main_LeafBlock94_SwitchLeaf95 == 1'd1))
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock94_SwitchLeaf95 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default13_i_79;
LEGUP_F_main_BB_LeafBlock99_90:
	if ((fsm_stall == 1'd0) && (1'd1 == 1'd1))
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
	else if ((fsm_stall == 1'd0) && (1'd1 == 1'd0))
		next_state = LEGUP_F_main_BB_LeafBlock99_sw_default31_i_crit_edge_91;
LEGUP_F_main_BB_LeafBlock99_sw_default31_i_crit_edge_91:
		next_state = LEGUP_F_main_BB_sw_default31_i_96;
LEGUP_F_main_BB_LeafBlock_24:
	if ((fsm_stall == 1'd0) && (main_LeafBlock_SwitchLeaf == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb118_i_34;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock_SwitchLeaf == 1'd0))
		next_state = LEGUP_F_main_BB_sw_default_i_35;
LEGUP_F_main_BB_NodeBlock101_89:
	if ((fsm_stall == 1'd0) && (main_NodeBlock101_Pivot102 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock99_90;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock101_Pivot102 == 1'd0))
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
LEGUP_F_main_BB_NodeBlock103_88:
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
LEGUP_F_main_BB_NodeBlock105_87:
	if ((fsm_stall == 1'd0) && (main_NodeBlock105_Pivot106 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock101_89;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock105_Pivot106 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock103_88;
LEGUP_F_main_BB_NodeBlock107_86:
	if ((fsm_stall == 1'd0) && (main_NodeBlock107_Pivot108 == 1'd1))
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock107_Pivot108 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock122_92;
LEGUP_F_main_BB_NodeBlock111_83:
	if ((fsm_stall == 1'd0) && (main_NodeBlock111_Pivot112 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock109_84;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock111_Pivot112 == 1'd0))
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
LEGUP_F_main_BB_NodeBlock113_82:
	if ((fsm_stall == 1'd0) && (main_NodeBlock113_Pivot114 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock107_86;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock113_Pivot114 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock111_83;
LEGUP_F_main_BB_NodeBlock115_81:
	if ((fsm_stall == 1'd0) && (main_NodeBlock115_Pivot116 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock105_87;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock115_Pivot116 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock113_82;
LEGUP_F_main_BB_NodeBlock11_17:
	if ((fsm_stall == 1'd0) && (main_NodeBlock11_Pivot12 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock3_21;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock11_Pivot12 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock9_18;
LEGUP_F_main_BB_NodeBlock122_92:
	if ((fsm_stall == 1'd0) && (main_NodeBlock122_Pivot123 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock118_94;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock122_Pivot123 == 1'd0))
		next_state = LEGUP_F_main_BB_LeafBlock120_93;
LEGUP_F_main_BB_NodeBlock127_130:
	if ((fsm_stall == 1'd0) && (main_NodeBlock127_Pivot128 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb1_i_132;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock127_Pivot128 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_bb5_i_133;
LEGUP_F_main_BB_NodeBlock129_129:
	if ((fsm_stall == 1'd0) && (main_NodeBlock129_Pivot130 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock125_131;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock129_Pivot130 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock127_130;
LEGUP_F_main_BB_NodeBlock131_128:
	if ((fsm_stall == 1'd0) && (main_NodeBlock131_Pivot132 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb13_i_135;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock131_Pivot132 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_bb17_i_136;
LEGUP_F_main_BB_NodeBlock133_127:
	if ((fsm_stall == 1'd0) && (main_NodeBlock133_Pivot134 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb9_i_134;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock133_Pivot134 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock131_128;
LEGUP_F_main_BB_NodeBlock135_126:
	if ((fsm_stall == 1'd0) && (main_NodeBlock135_Pivot136 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock129_129;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock135_Pivot136 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock133_127;
LEGUP_F_main_BB_NodeBlock137_125:
	if ((fsm_stall == 1'd0) && (main_NodeBlock137_Pivot138 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb31_i_138;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock137_Pivot138 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_bb37_i_139;
LEGUP_F_main_BB_NodeBlock139_124:
	if ((fsm_stall == 1'd0) && (main_NodeBlock139_Pivot140 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb22_i_137;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock139_Pivot140 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock137_125;
LEGUP_F_main_BB_NodeBlock141_123:
	if ((fsm_stall == 1'd0) && (main_NodeBlock141_Pivot142 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb49_i_141;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock141_Pivot142 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_bb54_i_142;
LEGUP_F_main_BB_NodeBlock143_122:
	if ((fsm_stall == 1'd0) && (main_NodeBlock143_Pivot144 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb42_i_140;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock143_Pivot144 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock141_123;
LEGUP_F_main_BB_NodeBlock145_121:
	if ((fsm_stall == 1'd0) && (main_NodeBlock145_Pivot146 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock139_124;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock145_Pivot146 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock143_122;
LEGUP_F_main_BB_NodeBlock147_120:
	if ((fsm_stall == 1'd0) && (main_NodeBlock147_Pivot148 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock135_126;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock147_Pivot148 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock145_121;
LEGUP_F_main_BB_NodeBlock149_119:
	if ((fsm_stall == 1'd0) && (main_NodeBlock149_Pivot150 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb65_i_144;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock149_Pivot150 == 1'd0))
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_NodeBlock151_118:
	if ((fsm_stall == 1'd0) && (main_NodeBlock151_Pivot152 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb60_i_143;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock151_Pivot152 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock149_119;
LEGUP_F_main_BB_NodeBlock153_117:
	if ((fsm_stall == 1'd0) && (main_NodeBlock153_Pivot154 == 1'd1))
		next_state = LEGUP_F_main_BB_alu_exit_154;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock153_Pivot154 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_bb83_i_147;
LEGUP_F_main_BB_NodeBlock155_116:
	if ((fsm_stall == 1'd0) && (main_NodeBlock155_Pivot156 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb73_i_146;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock155_Pivot156 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock153_117;
LEGUP_F_main_BB_NodeBlock157_115:
	if ((fsm_stall == 1'd0) && (main_NodeBlock157_Pivot158 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock151_118;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock157_Pivot158 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock155_116;
LEGUP_F_main_BB_NodeBlock161_113:
	if ((fsm_stall == 1'd0) && (main_NodeBlock161_Pivot162 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock159_114;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock161_Pivot162 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_bb106_i_150;
LEGUP_F_main_BB_NodeBlock163_112:
	if ((fsm_stall == 1'd0) && (main_NodeBlock163_Pivot164 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb88_i_148;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock163_Pivot164 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock161_113;
LEGUP_F_main_BB_NodeBlock167_110:
	if ((fsm_stall == 1'd0) && (main_NodeBlock167_Pivot168 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb124_i_152;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock167_Pivot168 == 1'd0))
		next_state = LEGUP_F_main_BB_LeafBlock165_111;
LEGUP_F_main_BB_NodeBlock169_109:
	if ((fsm_stall == 1'd0) && (main_NodeBlock169_Pivot170 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb115_i_151;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock169_Pivot170 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock167_110;
LEGUP_F_main_BB_NodeBlock171_108:
	if ((fsm_stall == 1'd0) && (main_NodeBlock171_Pivot172 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock163_112;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock171_Pivot172 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock169_109;
LEGUP_F_main_BB_NodeBlock173_107:
	if ((fsm_stall == 1'd0) && (main_NodeBlock173_Pivot174 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock157_115;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock173_Pivot174 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock171_108;
LEGUP_F_main_BB_NodeBlock175_106:
	if ((fsm_stall == 1'd0) && (main_NodeBlock175_Pivot176 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock147_120;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock175_Pivot176 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock173_107;
LEGUP_F_main_BB_NodeBlock22_39:
	if ((fsm_stall == 1'd0) && (main_NodeBlock22_Pivot23 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock18_41;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock22_Pivot23 == 1'd0))
		next_state = LEGUP_F_main_BB_LeafBlock20_40;
LEGUP_F_main_BB_NodeBlock24_38:
	if ((fsm_stall == 1'd0) && (main_NodeBlock24_Pivot25 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock16_42;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock24_Pivot25 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock22_39;
LEGUP_F_main_BB_NodeBlock31_50:
	if ((fsm_stall == 1'd0) && (main_NodeBlock31_Pivot32 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock27_52;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock31_Pivot32 == 1'd0))
		next_state = LEGUP_F_main_BB_LeafBlock29_51;
LEGUP_F_main_BB_NodeBlock39_46:
	if ((fsm_stall == 1'd0) && (main_while_body_Pivot14_reg == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock35_48;
	else if ((fsm_stall == 1'd0) && (main_while_body_Pivot14_reg == 1'd0))
		next_state = LEGUP_F_main_BB_LeafBlock37_47;
LEGUP_F_main_BB_NodeBlock41_45:
	if ((fsm_stall == 1'd0) && (main_NodeBlock41_Pivot42 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock33_49;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock41_Pivot42 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock39_46;
LEGUP_F_main_BB_NodeBlock43_44:
	if ((fsm_stall == 1'd0) && (main_NodeBlock43_Pivot44 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock31_50;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock43_Pivot44 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock41_45;
LEGUP_F_main_BB_NodeBlock50_68:
	if ((fsm_stall == 1'd0) && (main_NodeBlock50_Pivot51 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock46_70;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock50_Pivot51 == 1'd0))
		next_state = LEGUP_F_main_BB_LeafBlock48_69;
LEGUP_F_main_BB_NodeBlock56_65:
	if ((fsm_stall == 1'd0) && (main_NodeBlock56_Pivot57 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock52_67;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock56_Pivot57 == 1'd0))
		next_state = LEGUP_F_main_BB_LeafBlock54_66;
LEGUP_F_main_BB_NodeBlock58_64:
	if ((fsm_stall == 1'd0) && (main_NodeBlock58_Pivot59 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock50_68;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock58_Pivot59 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock56_65;
LEGUP_F_main_BB_NodeBlock64_61:
	if ((fsm_stall == 1'd0) && (main_while_body_Pivot14_reg == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock60_63;
	else if ((fsm_stall == 1'd0) && (main_while_body_Pivot14_reg == 1'd0))
		next_state = LEGUP_F_main_BB_LeafBlock62_62;
LEGUP_F_main_BB_NodeBlock72_57:
	if ((fsm_stall == 1'd0) && (main_NodeBlock72_Pivot73 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock68_59;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock72_Pivot73 == 1'd0))
		next_state = LEGUP_F_main_BB_LeafBlock70_58;
LEGUP_F_main_BB_NodeBlock74_56:
	if ((fsm_stall == 1'd0) && (main_NodeBlock74_Pivot75 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock66_60;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock74_Pivot75 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock72_57;
LEGUP_F_main_BB_NodeBlock76_55:
	if ((fsm_stall == 1'd0) && (main_NodeBlock76_Pivot77 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock64_61;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock76_Pivot77 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock74_56;
LEGUP_F_main_BB_NodeBlock78_54:
	if ((fsm_stall == 1'd0) && (main_NodeBlock78_Pivot79 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock58_64;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock78_Pivot79 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock76_55;
LEGUP_F_main_BB_NodeBlock87_72:
	if ((fsm_stall == 1'd0) && (main_NodeBlock87_Pivot88 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock83_74;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock87_Pivot88 == 1'd0))
		next_state = LEGUP_F_main_BB_LeafBlock85_73;
LEGUP_F_main_BB_NodeBlock89_71:
	if ((fsm_stall == 1'd0) && (main_NodeBlock89_Pivot90 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock81_75;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock89_Pivot90 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock87_72;
LEGUP_F_main_BB_NodeBlock96_76:
	if ((fsm_stall == 1'd0) && (main_NodeBlock96_Pivot97 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock92_78;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock96_Pivot97 == 1'd0))
		next_state = LEGUP_F_main_BB_LeafBlock94_77;
LEGUP_F_main_BB_NodeBlock9_18:
	if ((fsm_stall == 1'd0) && (main_NodeBlock9_Pivot10 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock5_20;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock9_Pivot10 == 1'd0))
		next_state = LEGUP_F_main_BB_LeafBlock7_19;
LEGUP_F_main_BB_NodeBlock_22:
	if ((fsm_stall == 1'd0) && (main_NodeBlock_Pivot == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock_24;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock_Pivot == 1'd0))
		next_state = LEGUP_F_main_BB_LeafBlock1_23;
LEGUP_F_main_BB_addressCalculator_exit_172:
	if ((fsm_stall == 1'd0) && (main_addressCalculator_exit_or_cond == 1'd1))
		next_state = LEGUP_F_main_BB_if_end61_while_body_crit_edge_173;
	else if ((fsm_stall == 1'd0) && (main_addressCalculator_exit_or_cond == 1'd0))
		next_state = LEGUP_F_main_BB_while_end_175;
LEGUP_F_main_BB_aluDecode_exit_102:
		next_state = LEGUP_F_main_BB_aluDecode_exit_103;
LEGUP_F_main_BB_aluDecode_exit_103:
	if ((fsm_stall == 1'd0) && (main_aluDecode_exit_tobool_reg == 1'd1))
		next_state = LEGUP_F_main_BB_if_else_104;
	else if ((fsm_stall == 1'd0) && (main_aluDecode_exit_tobool_reg == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock175_106;
LEGUP_F_main_BB_alu_exit_154:
	if ((fsm_stall == 1'd0) && (main_alu_exit_tobool34 == 1'd1))
		next_state = LEGUP_F_main_BB_if_end42_158;
	else if ((fsm_stall == 1'd0) && (main_alu_exit_tobool34 == 1'd0))
		next_state = LEGUP_F_main_BB_if_then38_155;
LEGUP_F_main_BB_if_else131_i_37:
		next_state = LEGUP_F_main_BB_NodeBlock24_38;
LEGUP_F_main_BB_if_else15_i_170:
		next_state = LEGUP_F_main_BB_addressCalculator_exit_172;
LEGUP_F_main_BB_if_else18_i_171:
		next_state = LEGUP_F_main_BB_addressCalculator_exit_172;
LEGUP_F_main_BB_if_else51_162:
	if ((fsm_stall == 1'd0) && (main_if_else51_tobool52 == 1'd1))
		next_state = LEGUP_F_main_BB_if_end61_165;
	else if ((fsm_stall == 1'd0) && (main_if_else51_tobool52 == 1'd0))
		next_state = LEGUP_F_main_BB_if_then56_163;
LEGUP_F_main_BB_if_else62_i_30:
		next_state = LEGUP_F_main_BB_sw_default148_i_53;
LEGUP_F_main_BB_if_else_104:
		next_state = LEGUP_F_main_BB_if_else_105;
LEGUP_F_main_BB_if_else_105:
		next_state = LEGUP_F_main_BB_NodeBlock175_106;
LEGUP_F_main_BB_if_else_i2_168:
	if ((fsm_stall == 1'd0) && (main_if_end61_tobool66_reg == 1'd1))
		next_state = LEGUP_F_main_BB_if_else15_i_170;
	else if ((fsm_stall == 1'd0) && (main_if_end61_tobool66_reg == 1'd0))
		next_state = LEGUP_F_main_BB_if_then13_i_169;
LEGUP_F_main_BB_if_else_i_27:
		next_state = LEGUP_F_main_BB_sw_default148_i_53;
LEGUP_F_main_BB_if_end42_158:
	if ((fsm_stall == 1'd0) && (main_if_end42_tobool43 == 1'd1))
		next_state = LEGUP_F_main_BB_if_else51_162;
	else if ((fsm_stall == 1'd0) && (main_if_end42_tobool43 == 1'd0))
		next_state = LEGUP_F_main_BB_if_then47_159;
LEGUP_F_main_BB_if_end61_165:
	if ((fsm_stall == 1'd0) && (main_if_end61_tobool63 == 1'd1))
		next_state = LEGUP_F_main_BB_if_else18_i_171;
	else if ((fsm_stall == 1'd0) && (main_if_end61_tobool63 == 1'd0))
		next_state = LEGUP_F_main_BB_if_then_i1_166;
LEGUP_F_main_BB_if_end61_while_body_crit_edge_173:
		next_state = LEGUP_F_main_BB_if_end61_while_body_crit_edge_174;
LEGUP_F_main_BB_if_end61_while_body_crit_edge_174:
		next_state = LEGUP_F_main_BB_while_body_15;
LEGUP_F_main_BB_if_then126_i_36:
		next_state = LEGUP_F_main_BB_NodeBlock24_38;
LEGUP_F_main_BB_if_then13_i_169:
		next_state = LEGUP_F_main_BB_addressCalculator_exit_172;
LEGUP_F_main_BB_if_then38_155:
		next_state = LEGUP_F_main_BB_if_then38_156;
LEGUP_F_main_BB_if_then38_156:
		next_state = LEGUP_F_main_BB_if_then38_157;
LEGUP_F_main_BB_if_then38_157:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_if_then44_i_29:
		next_state = LEGUP_F_main_BB_NodeBlock24_38;
LEGUP_F_main_BB_if_then47_159:
		next_state = LEGUP_F_main_BB_if_then47_160;
LEGUP_F_main_BB_if_then47_160:
		next_state = LEGUP_F_main_BB_if_then47_161;
LEGUP_F_main_BB_if_then47_161:
		next_state = LEGUP_F_main_BB_if_end61_165;
LEGUP_F_main_BB_if_then56_163:
		next_state = LEGUP_F_main_BB_if_then56_164;
LEGUP_F_main_BB_if_then56_164:
		next_state = LEGUP_F_main_BB_if_end61_165;
LEGUP_F_main_BB_if_then88_i_32:
		next_state = LEGUP_F_main_BB_NodeBlock24_38;
LEGUP_F_main_BB_if_then8_i_167:
		next_state = LEGUP_F_main_BB_addressCalculator_exit_172;
LEGUP_F_main_BB_if_then_i1_166:
	if ((fsm_stall == 1'd0) && (main_if_then_i1_tobool65 == 1'd1))
		next_state = LEGUP_F_main_BB_if_else_i2_168;
	else if ((fsm_stall == 1'd0) && (main_if_then_i1_tobool65 == 1'd0))
		next_state = LEGUP_F_main_BB_if_then8_i_167;
LEGUP_F_main_BB_if_then_i_26:
		next_state = LEGUP_F_main_BB_NodeBlock24_38;
LEGUP_F_main_BB_legup_memset_4_exit_10:
		next_state = LEGUP_F_main_BB_legup_memset_4_exit_11;
LEGUP_F_main_BB_legup_memset_4_exit_11:
		next_state = LEGUP_F_main_BB_legup_memset_4_exit_12;
LEGUP_F_main_BB_legup_memset_4_exit_12:
		next_state = LEGUP_F_main_BB_legup_memset_4_exit_13;
LEGUP_F_main_BB_legup_memset_4_exit_13:
		next_state = LEGUP_F_main_BB_legup_memset_4_exit_14;
LEGUP_F_main_BB_legup_memset_4_exit_14:
		next_state = LEGUP_F_main_BB_while_body_15;
LEGUP_F_main_BB_legup_memset_4_exit_4:
		next_state = LEGUP_F_main_BB_legup_memset_4_exit_5;
LEGUP_F_main_BB_legup_memset_4_exit_5:
		next_state = LEGUP_F_main_BB_legup_memset_4_exit_6;
LEGUP_F_main_BB_legup_memset_4_exit_6:
		next_state = LEGUP_F_main_BB_legup_memset_4_exit_7;
LEGUP_F_main_BB_legup_memset_4_exit_7:
		next_state = LEGUP_F_main_BB_legup_memset_4_exit_8;
LEGUP_F_main_BB_legup_memset_4_exit_8:
		next_state = LEGUP_F_main_BB_legup_memset_4_exit_9;
LEGUP_F_main_BB_legup_memset_4_exit_9:
		next_state = LEGUP_F_main_BB_legup_memset_4_exit_10;
LEGUP_F_main_BB_sw_bb106_i_150:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb115_i_151:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb118_i_34:
		next_state = LEGUP_F_main_BB_NodeBlock24_38;
LEGUP_F_main_BB_sw_bb124_i_152:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb133_i_153:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb13_i_135:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb17_i_136:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb1_i_132:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb22_i_137:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb31_i_138:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb37_i_139:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb40_i_28:
	if ((fsm_stall == 1'd0) && (main_sw_bb40_i_cmp43_i == 1'd1))
		next_state = LEGUP_F_main_BB_if_then44_i_29;
	else if ((fsm_stall == 1'd0) && (main_sw_bb40_i_cmp43_i == 1'd0))
		next_state = LEGUP_F_main_BB_if_else62_i_30;
LEGUP_F_main_BB_sw_bb42_i_140:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb49_i_141:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb54_i_142:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb5_i_133:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb60_i_143:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb65_i_144:
		next_state = LEGUP_F_main_BB_sw_bb65_i_145;
LEGUP_F_main_BB_sw_bb65_i_145:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb73_i_146:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb83_i_147:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb84_i_31:
	if ((fsm_stall == 1'd0) && (main_sw_bb84_i_cmp87_i == 1'd1))
		next_state = LEGUP_F_main_BB_if_then88_i_32;
	else if ((fsm_stall == 1'd0) && (main_sw_bb84_i_cmp87_i == 1'd0))
		next_state = LEGUP_F_main_BB_sw_epilog_thread242_i_33;
LEGUP_F_main_BB_sw_bb88_i_148:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb97_i_149:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb9_i_134:
		next_state = LEGUP_F_main_BB_if_end42_158;
LEGUP_F_main_BB_sw_bb_i_25:
	if ((fsm_stall == 1'd0) && (main_sw_bb_i_cmp_i == 1'd1))
		next_state = LEGUP_F_main_BB_if_then_i_26;
	else if ((fsm_stall == 1'd0) && (main_sw_bb_i_cmp_i == 1'd0))
		next_state = LEGUP_F_main_BB_if_else_i_27;
LEGUP_F_main_BB_sw_default13_i_79:
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
LEGUP_F_main_BB_sw_default142_i_43:
		next_state = LEGUP_F_main_BB_NodeBlock43_44;
LEGUP_F_main_BB_sw_default148_i_53:
		next_state = LEGUP_F_main_BB_NodeBlock78_54;
LEGUP_F_main_BB_sw_default16_i_80:
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
LEGUP_F_main_BB_sw_default29_i_95:
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
LEGUP_F_main_BB_sw_default31_i_96:
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
LEGUP_F_main_BB_sw_default48_i_97:
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
LEGUP_F_main_BB_sw_default_i_35:
	if ((fsm_stall == 1'd0) && (main_while_body_bit_select16_reg == 1'd1))
		next_state = LEGUP_F_main_BB_if_then126_i_36;
	else if ((fsm_stall == 1'd0) && (main_while_body_bit_select16_reg == 1'd0))
		next_state = LEGUP_F_main_BB_if_else131_i_37;
LEGUP_F_main_BB_sw_epilog_thread242_i_33:
		next_state = LEGUP_F_main_BB_sw_default142_i_43;
LEGUP_F_main_BB_switch_lookup54_i_100:
		next_state = LEGUP_F_main_BB_switch_lookup54_i_101;
LEGUP_F_main_BB_switch_lookup54_i_101:
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
LEGUP_F_main_BB_switch_lookup_i_98:
		next_state = LEGUP_F_main_BB_switch_lookup_i_99;
LEGUP_F_main_BB_switch_lookup_i_99:
		next_state = LEGUP_F_main_BB_aluDecode_exit_102;
LEGUP_F_main_BB_while_body_15:
		next_state = LEGUP_F_main_BB_while_body_16;
LEGUP_F_main_BB_while_body_16:
	if ((fsm_stall == 1'd0) && (main_while_body_Pivot14_reg == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock_22;
	else if ((fsm_stall == 1'd0) && (main_while_body_Pivot14_reg == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock11_17;
LEGUP_F_main_BB_while_body_i_2:
		next_state = LEGUP_F_main_BB_while_body_i_3;
LEGUP_F_main_BB_while_body_i_3:
	if ((fsm_stall == 1'd0) && (main_while_body_i_exitcond1_reg == 1'd1))
		next_state = LEGUP_F_main_BB_legup_memset_4_exit_4;
	else if ((fsm_stall == 1'd0) && (main_while_body_i_exitcond1_reg == 1'd0))
		next_state = LEGUP_F_main_BB_while_body_i_2;
LEGUP_F_main_BB_while_body_lr_ph_1:
		next_state = LEGUP_F_main_BB_while_body_i_2;
LEGUP_F_main_BB_while_end_175:
		next_state = LEGUP_F_main_BB_while_end_176;
LEGUP_F_main_BB_while_end_176:
		next_state = LEGUP_0;
default:
	next_state = cur_state;
endcase

end
assign fsm_stall = 1'd0;
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_while_body_lr_ph_1) & (fsm_stall == 1'd0))) begin
		main_while_body_i_indvar = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_while_body_i_3) & (fsm_stall == 1'd0)) & (main_while_body_i_exitcond1_reg == 1'd0))) */ begin
		main_while_body_i_indvar = main_while_body_i_0_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_while_body_lr_ph_1) & (fsm_stall == 1'd0))) begin
		main_while_body_i_indvar_reg <= main_while_body_i_indvar;
	end
	if ((((cur_state == LEGUP_F_main_BB_while_body_i_3) & (fsm_stall == 1'd0)) & (main_while_body_i_exitcond1_reg == 1'd0))) begin
		main_while_body_i_indvar_reg <= main_while_body_i_indvar;
	end
end
always @(*) begin
		main_while_body_i_s_010_i = (1'd0 + (4 * {26'd0,main_while_body_i_indvar_reg}));
end
always @(*) begin
		main_while_body_i_0 = ({1'd0,main_while_body_i_indvar_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_i_2)) begin
		main_while_body_i_0_reg <= main_while_body_i_0;
	end
end
always @(*) begin
		main_while_body_i_exitcond1 = (main_while_body_i_0 == 32'd32);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_i_2)) begin
		main_while_body_i_exitcond1_reg <= main_while_body_i_exitcond1;
	end
end
assign main_legup_memset_4_exit_arrayidx = 1'd0;
assign main_legup_memset_4_exit_arrayidx1 = (1'd0 + (4 * 32'd4));
assign main_legup_memset_4_exit_arrayidx2 = (1'd0 + (4 * 32'd8));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx2_reg <= main_legup_memset_4_exit_arrayidx2;
	end
end
assign main_legup_memset_4_exit_arrayidx3 = (1'd0 + (4 * 32'd12));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx3_reg <= main_legup_memset_4_exit_arrayidx3;
	end
end
assign main_legup_memset_4_exit_arrayidx4 = (1'd0 + (4 * 32'd16));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx4_reg <= main_legup_memset_4_exit_arrayidx4;
	end
end
assign main_legup_memset_4_exit_arrayidx5 = (1'd0 + (4 * 32'd20));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx5_reg <= main_legup_memset_4_exit_arrayidx5;
	end
end
assign main_legup_memset_4_exit_arrayidx6 = (1'd0 + (4 * 32'd24));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx6_reg <= main_legup_memset_4_exit_arrayidx6;
	end
end
assign main_legup_memset_4_exit_arrayidx7 = (1'd0 + (4 * 32'd28));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx7_reg <= main_legup_memset_4_exit_arrayidx7;
	end
end
assign main_legup_memset_4_exit_arrayidx8 = (1'd0 + (4 * 32'd32));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx8_reg <= main_legup_memset_4_exit_arrayidx8;
	end
end
assign main_legup_memset_4_exit_arrayidx9 = (1'd0 + (4 * 32'd36));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx9_reg <= main_legup_memset_4_exit_arrayidx9;
	end
end
assign main_legup_memset_4_exit_arrayidx10 = (1'd0 + (4 * 32'd40));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx10_reg <= main_legup_memset_4_exit_arrayidx10;
	end
end
assign main_legup_memset_4_exit_arrayidx11 = (1'd0 + (4 * 32'd44));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx11_reg <= main_legup_memset_4_exit_arrayidx11;
	end
end
assign main_legup_memset_4_exit_arrayidx12 = (1'd0 + (4 * 32'd48));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx12_reg <= main_legup_memset_4_exit_arrayidx12;
	end
end
assign main_legup_memset_4_exit_arrayidx13 = (1'd0 + (4 * 32'd52));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx13_reg <= main_legup_memset_4_exit_arrayidx13;
	end
end
assign main_legup_memset_4_exit_arrayidx14 = (1'd0 + (4 * 32'd56));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx14_reg <= main_legup_memset_4_exit_arrayidx14;
	end
end
assign main_legup_memset_4_exit_arrayidx15 = (1'd0 + (4 * 32'd60));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx15_reg <= main_legup_memset_4_exit_arrayidx15;
	end
end
assign main_legup_memset_4_exit_arrayidx16 = (1'd0 + (4 * 32'd64));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx16_reg <= main_legup_memset_4_exit_arrayidx16;
	end
end
assign main_legup_memset_4_exit_arrayidx17 = (1'd0 + (4 * 32'd68));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx17_reg <= main_legup_memset_4_exit_arrayidx17;
	end
end
assign main_legup_memset_4_exit_arrayidx18 = (1'd0 + (4 * 32'd72));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx18_reg <= main_legup_memset_4_exit_arrayidx18;
	end
end
assign main_legup_memset_4_exit_arrayidx19 = (1'd0 + (4 * 32'd76));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx19_reg <= main_legup_memset_4_exit_arrayidx19;
	end
end
assign main_legup_memset_4_exit_arrayidx22 = 1'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_legup_memset_4_exit_arrayidx22_reg <= main_legup_memset_4_exit_arrayidx22;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_14) & (fsm_stall == 1'd0))) begin
		main_while_body_1 = 32'd536871187;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_if_end61_while_body_crit_edge_174) & (fsm_stall == 1'd0))) */ begin
		main_while_body_1 = main_if_end61_while_body_crit_edge_pre100;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_14) & (fsm_stall == 1'd0))) begin
		main_while_body_1_reg <= main_while_body_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end61_while_body_crit_edge_174) & (fsm_stall == 1'd0))) begin
		main_while_body_1_reg <= main_while_body_1;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_14) & (fsm_stall == 1'd0))) begin
		main_while_body_nextInst_099 = 32'd0;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_if_end61_while_body_crit_edge_174) & (fsm_stall == 1'd0))) */ begin
		main_while_body_nextInst_099 = main_addressCalculator_exit_newPc_0_i_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_14) & (fsm_stall == 1'd0))) begin
		main_while_body_nextInst_099_reg <= main_while_body_nextInst_099;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end61_while_body_crit_edge_174) & (fsm_stall == 1'd0))) begin
		main_while_body_nextInst_099_reg <= main_while_body_nextInst_099;
	end
end
always @(*) begin
		main_while_body_bit_select44 = main_while_body_1_reg[19:15];
end
always @(*) begin
		main_while_body_bit_select42 = main_while_body_1_reg[24:20];
end
always @(*) begin
		main_while_body_bit_select39 = main_while_body_1_reg[14:12];
end
always @(*) begin
		main_while_body_bit_select37 = main_while_body_1_reg[6:0];
end
always @(*) begin
		main_while_body_bit_select32 = main_while_body_1_reg[30:21];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_bit_select32_reg <= main_while_body_bit_select32;
	end
end
always @(*) begin
		main_while_body_bit_select30 = main_while_body_1_reg[24:21];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_bit_select30_reg <= main_while_body_bit_select30;
	end
end
always @(*) begin
		main_while_body_bit_select29 = main_while_body_1_reg[20];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_bit_select29_reg <= main_while_body_bit_select29;
	end
end
always @(*) begin
		main_while_body_bit_select28 = main_while_body_1_reg[19:12];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_bit_select28_reg <= main_while_body_bit_select28;
	end
end
always @(*) begin
		main_while_body_bit_select25 = main_while_body_1_reg[7];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_bit_select25_reg <= main_while_body_bit_select25;
	end
end
always @(*) begin
		main_while_body_bit_select24 = main_while_body_1_reg[11:8];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_bit_select24_reg <= main_while_body_bit_select24;
	end
end
always @(*) begin
		main_while_body_bit_select23 = main_while_body_1_reg[29:25];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_bit_select23_reg <= main_while_body_bit_select23;
	end
end
always @(*) begin
		main_while_body_bit_select21 = main_while_body_1_reg[11:7];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_bit_select21_reg <= main_while_body_bit_select21;
	end
end
always @(*) begin
		main_while_body_bit_select20 = main_while_body_1_reg[30:25];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_bit_select20_reg <= main_while_body_bit_select20;
	end
end
always @(*) begin
		main_while_body_bit_select17 = main_while_body_1_reg[31:12];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_bit_select17_reg <= main_while_body_bit_select17;
	end
end
always @(*) begin
		main_while_body_bit_select16 = main_while_body_1_reg[31];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_bit_select16_reg <= main_while_body_bit_select16;
	end
end
always @(*) begin
		main_while_body_bit_select13 = main_while_body_1_reg[30:20];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_bit_select13_reg <= main_while_body_bit_select13;
	end
end
always @(*) begin
		main_while_body_bit_concat45 = {main_while_body_bit_concat45_bit_select_operand_0[26:0], main_while_body_bit_select44[4:0]};
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_bit_concat45_reg <= main_while_body_bit_concat45;
	end
end
always @(*) begin
		main_while_body_bit_concat43 = {main_while_body_bit_concat43_bit_select_operand_0[26:0], main_while_body_bit_select42[4:0]};
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_bit_concat43_reg <= main_while_body_bit_concat43;
	end
end
always @(*) begin
		main_while_body_bit_concat41 = {main_while_body_bit_concat41_bit_select_operand_0[26:0], main_while_body_bit_select21[4:0]};
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_bit_concat41_reg <= main_while_body_bit_concat41;
	end
end
always @(*) begin
		main_while_body_shr6_i = ($signed(main_while_body_1_reg) >>> 32'd25);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_shr6_i_reg <= main_while_body_shr6_i;
	end
end
always @(*) begin
		main_while_body_bit_concat40 = {main_while_body_bit_concat40_bit_select_operand_0[28:0], main_while_body_bit_select39[2:0]};
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_bit_concat40_reg <= main_while_body_bit_concat40;
	end
end
always @(*) begin
		main_while_body_bit_concat38 = {main_while_body_bit_concat38_bit_select_operand_0[24:0], main_while_body_bit_select37[6:0]};
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_bit_concat38_reg <= main_while_body_bit_concat38;
	end
end
always @(*) begin
		main_while_body_Pivot14 = (main_while_body_bit_concat38 < 32'd55);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_Pivot14_reg <= main_while_body_Pivot14;
	end
end
always @(*) begin
		main_NodeBlock11_Pivot12 = (main_while_body_bit_concat38_reg < 32'd99);
end
always @(*) begin
		main_NodeBlock9_Pivot10 = (main_while_body_bit_concat38_reg < 32'd111);
end
always @(*) begin
		main_LeafBlock7_SwitchLeaf8 = (main_while_body_bit_concat38_reg == 32'd111);
end
always @(*) begin
		main_LeafBlock5_SwitchLeaf6 = (main_while_body_bit_concat38_reg == 32'd99);
end
always @(*) begin
		main_LeafBlock3_SwitchLeaf4 = (main_while_body_bit_concat38_reg == 32'd55);
end
always @(*) begin
		main_NodeBlock_Pivot = (main_while_body_bit_concat38_reg < 32'd35);
end
always @(*) begin
		main_LeafBlock1_SwitchLeaf2 = (main_while_body_bit_concat38_reg == 32'd35);
end
always @(*) begin
		main_LeafBlock_SwitchLeaf = (main_while_body_bit_concat38_reg == 32'd23);
end
always @(*) begin
		main_sw_bb_i_shr13_i = ($signed(main_while_body_1_reg) >>> 32'd31);
end
always @(*) begin
		main_sw_bb_i_bit_select34 = main_sw_bb_i_shr13_i[0];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_sw_bb_i_25)) begin
		main_sw_bb_i_bit_select34_reg <= main_sw_bb_i_bit_select34;
	end
end
always @(*) begin
		main_sw_bb_i_cmp_i = ($signed(main_sw_bb_i_shr13_i) == $signed(-32'd1));
end
always @(*) begin
		main_if_then_i_bit_concat36 = {{{main_if_then_i_bit_concat36_bit_select_operand_0[20:0], main_while_body_bit_select20_reg[5:0]}, main_while_body_bit_select24_reg[3:0]}, main_if_then_i_bit_concat36_bit_select_operand_6};
end
always @(*) begin
		main_if_else_i_bit_concat35 = {{{{{{main_sw_bb_i_bit_select34_reg, main_if_else_i_bit_concat35_bit_select_operand_2[17:0]}, main_while_body_bit_select25_reg}, main_if_else_i_bit_concat35_bit_select_operand_6}, main_while_body_bit_select20_reg[5:0]}, main_while_body_bit_select24_reg[3:0]}, main_if_else_i_bit_concat35_bit_select_operand_12};
end
always @(*) begin
		main_sw_bb40_i_shr42_i = ($signed(main_while_body_1_reg) >>> 32'd31);
end
always @(*) begin
		main_sw_bb40_i_bit_select27 = main_sw_bb40_i_shr42_i[0];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_sw_bb40_i_28)) begin
		main_sw_bb40_i_bit_select27_reg <= main_sw_bb40_i_bit_select27;
	end
end
always @(*) begin
		main_sw_bb40_i_cmp43_i = ($signed(main_sw_bb40_i_shr42_i) == $signed(-32'd1));
end
always @(*) begin
		main_if_then44_i_bit_concat33 = {{{{main_if_then44_i_bit_concat33_bit_select_operand_0[11:0], main_while_body_bit_select28_reg[7:0]}, main_while_body_bit_select29_reg}, main_while_body_bit_select32_reg[9:0]}, main_if_then44_i_bit_concat33_bit_select_operand_8};
end
always @(*) begin
		main_if_else62_i_bit_concat31 = {{{{{{main_sw_bb40_i_bit_select27_reg, main_if_else62_i_bit_concat31_bit_select_operand_2[10:0]}, main_while_body_bit_select28_reg[7:0]}, main_while_body_bit_select29_reg}, main_while_body_bit_select20_reg[5:0]}, main_while_body_bit_select30_reg[3:0]}, main_if_else62_i_bit_concat31_bit_select_operand_12};
end
always @(*) begin
		main_sw_bb84_i_shr86_i = ($signed(main_while_body_1_reg) >>> 32'd31);
end
always @(*) begin
		main_sw_bb84_i_bit_select19 = main_sw_bb84_i_shr86_i[0];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_sw_bb84_i_31)) begin
		main_sw_bb84_i_bit_select19_reg <= main_sw_bb84_i_bit_select19;
	end
end
always @(*) begin
		main_sw_bb84_i_cmp87_i = ($signed(main_sw_bb84_i_shr86_i) == $signed(-32'd1));
end
always @(*) begin
		main_if_then88_i_bit_concat26 = {{{{main_if_then88_i_bit_concat26_bit_select_operand_0[20:0], main_while_body_bit_select23_reg[4:0]}, main_if_then88_i_bit_concat26_bit_select_operand_4}, main_while_body_bit_select24_reg[3:0]}, main_while_body_bit_select25_reg};
end
always @(*) begin
		main_sw_epilog_thread242_i_bit_concat22 = {{{{main_sw_bb84_i_bit_select19_reg, main_sw_epilog_thread242_i_bit_concat22_bit_select_operand_2[18:0]}, main_while_body_bit_select20_reg[5:0]}, main_sw_epilog_thread242_i_bit_concat22_bit_select_operand_6}, main_while_body_bit_select21_reg[4:0]};
end
always @(*) begin
		main_sw_bb118_i_bit_concat18 = {main_while_body_bit_select17_reg[19:0], main_sw_bb118_i_bit_concat18_bit_select_operand_2[11:0]};
end
always @(*) begin
		main_if_then126_i_bit_concat15 = {main_if_then126_i_bit_concat15_bit_select_operand_0[20:0], main_while_body_bit_select13_reg[10:0]};
end
always @(*) begin
		main_if_else131_i_bit_concat14 = {main_if_else131_i_bit_concat14_bit_select_operand_0[20:0], main_while_body_bit_select13_reg[10:0]};
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_if_then_i_26) & (fsm_stall == 1'd0))) begin
		main_NodeBlock24_results_sroa_14_0_i = main_if_then_i_bit_concat36;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_then44_i_29) & (fsm_stall == 1'd0))) begin
		main_NodeBlock24_results_sroa_14_0_i = main_if_then44_i_bit_concat33;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_then88_i_32) & (fsm_stall == 1'd0))) begin
		main_NodeBlock24_results_sroa_14_0_i = main_if_then88_i_bit_concat26;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb118_i_34) & (fsm_stall == 1'd0))) begin
		main_NodeBlock24_results_sroa_14_0_i = main_sw_bb118_i_bit_concat18;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_then126_i_36) & (fsm_stall == 1'd0))) begin
		main_NodeBlock24_results_sroa_14_0_i = main_if_then126_i_bit_concat15;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_if_else131_i_37) & (fsm_stall == 1'd0))) */ begin
		main_NodeBlock24_results_sroa_14_0_i = main_if_else131_i_bit_concat14;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_if_then_i_26) & (fsm_stall == 1'd0))) begin
		main_NodeBlock24_results_sroa_14_0_i_reg <= main_NodeBlock24_results_sroa_14_0_i;
	end
	if (((cur_state == LEGUP_F_main_BB_if_then44_i_29) & (fsm_stall == 1'd0))) begin
		main_NodeBlock24_results_sroa_14_0_i_reg <= main_NodeBlock24_results_sroa_14_0_i;
	end
	if (((cur_state == LEGUP_F_main_BB_if_then88_i_32) & (fsm_stall == 1'd0))) begin
		main_NodeBlock24_results_sroa_14_0_i_reg <= main_NodeBlock24_results_sroa_14_0_i;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb118_i_34) & (fsm_stall == 1'd0))) begin
		main_NodeBlock24_results_sroa_14_0_i_reg <= main_NodeBlock24_results_sroa_14_0_i;
	end
	if (((cur_state == LEGUP_F_main_BB_if_then126_i_36) & (fsm_stall == 1'd0))) begin
		main_NodeBlock24_results_sroa_14_0_i_reg <= main_NodeBlock24_results_sroa_14_0_i;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else131_i_37) & (fsm_stall == 1'd0))) begin
		main_NodeBlock24_results_sroa_14_0_i_reg <= main_NodeBlock24_results_sroa_14_0_i;
	end
end
always @(*) begin
		main_NodeBlock24_Pivot25 = (main_while_body_bit_concat38_reg < 32'd103);
end
always @(*) begin
		main_NodeBlock22_Pivot23 = (main_while_body_bit_concat38_reg < 32'd111);
end
always @(*) begin
		main_LeafBlock20_SwitchLeaf21 = (main_while_body_bit_concat38_reg == 32'd111);
end
always @(*) begin
		main_LeafBlock18_SwitchLeaf19 = (main_while_body_bit_concat38_reg == 32'd103);
end
always @(*) begin
		main_LeafBlock16_SwitchLeaf17 = (main_while_body_bit_concat38_reg == 32'd99);
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_sw_epilog_thread242_i_33) & (fsm_stall == 1'd0))) begin
		main_sw_default142_i_results_sroa_14_0243_i = main_sw_epilog_thread242_i_bit_concat22;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock20_40) & (fsm_stall == 1'd0)) & (main_LeafBlock20_SwitchLeaf21 == 1'd0))) begin
		main_sw_default142_i_results_sroa_14_0243_i = main_NodeBlock24_results_sroa_14_0_i_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock18_41) & (fsm_stall == 1'd0)) & (main_LeafBlock18_SwitchLeaf19 == 1'd0))) begin
		main_sw_default142_i_results_sroa_14_0243_i = main_NodeBlock24_results_sroa_14_0_i_reg;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_LeafBlock16_42) & (fsm_stall == 1'd0)) & (main_LeafBlock16_SwitchLeaf17 == 1'd0))) */ begin
		main_sw_default142_i_results_sroa_14_0243_i = main_NodeBlock24_results_sroa_14_0_i_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_sw_epilog_thread242_i_33) & (fsm_stall == 1'd0))) begin
		main_sw_default142_i_results_sroa_14_0243_i_reg <= main_sw_default142_i_results_sroa_14_0243_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock20_40) & (fsm_stall == 1'd0)) & (main_LeafBlock20_SwitchLeaf21 == 1'd0))) begin
		main_sw_default142_i_results_sroa_14_0243_i_reg <= main_sw_default142_i_results_sroa_14_0243_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock18_41) & (fsm_stall == 1'd0)) & (main_LeafBlock18_SwitchLeaf19 == 1'd0))) begin
		main_sw_default142_i_results_sroa_14_0243_i_reg <= main_sw_default142_i_results_sroa_14_0243_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock16_42) & (fsm_stall == 1'd0)) & (main_LeafBlock16_SwitchLeaf17 == 1'd0))) begin
		main_sw_default142_i_results_sroa_14_0243_i_reg <= main_sw_default142_i_results_sroa_14_0243_i;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock20_40) & (fsm_stall == 1'd0)) & (main_LeafBlock20_SwitchLeaf21 == 1'd1))) begin
		main_NodeBlock43_results_sroa_14_0241_i = main_NodeBlock24_results_sroa_14_0_i_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock16_42) & (fsm_stall == 1'd0)) & (main_LeafBlock16_SwitchLeaf17 == 1'd1))) begin
		main_NodeBlock43_results_sroa_14_0241_i = main_NodeBlock24_results_sroa_14_0_i_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_sw_default142_i_43) & (fsm_stall == 1'd0))) */ begin
		main_NodeBlock43_results_sroa_14_0241_i = main_sw_default142_i_results_sroa_14_0243_i_reg;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock20_40) & (fsm_stall == 1'd0)) & (main_LeafBlock20_SwitchLeaf21 == 1'd1))) begin
		main_NodeBlock43_results_sroa_14_0241_i_reg <= main_NodeBlock43_results_sroa_14_0241_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock16_42) & (fsm_stall == 1'd0)) & (main_LeafBlock16_SwitchLeaf17 == 1'd1))) begin
		main_NodeBlock43_results_sroa_14_0241_i_reg <= main_NodeBlock43_results_sroa_14_0241_i;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default142_i_43) & (fsm_stall == 1'd0))) begin
		main_NodeBlock43_results_sroa_14_0241_i_reg <= main_NodeBlock43_results_sroa_14_0241_i;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock20_40) & (fsm_stall == 1'd0)) & (main_LeafBlock20_SwitchLeaf21 == 1'd1))) begin
		main_NodeBlock43_results_sroa_23_0_i = 8'd1;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock16_42) & (fsm_stall == 1'd0)) & (main_LeafBlock16_SwitchLeaf17 == 1'd1))) begin
		main_NodeBlock43_results_sroa_23_0_i = 8'd1;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_sw_default142_i_43) & (fsm_stall == 1'd0))) */ begin
		main_NodeBlock43_results_sroa_23_0_i = 8'd0;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock20_40) & (fsm_stall == 1'd0)) & (main_LeafBlock20_SwitchLeaf21 == 1'd1))) begin
		main_NodeBlock43_results_sroa_23_0_i_reg <= main_NodeBlock43_results_sroa_23_0_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock16_42) & (fsm_stall == 1'd0)) & (main_LeafBlock16_SwitchLeaf17 == 1'd1))) begin
		main_NodeBlock43_results_sroa_23_0_i_reg <= main_NodeBlock43_results_sroa_23_0_i;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default142_i_43) & (fsm_stall == 1'd0))) begin
		main_NodeBlock43_results_sroa_23_0_i_reg <= main_NodeBlock43_results_sroa_23_0_i;
	end
end
always @(*) begin
		main_NodeBlock43_Pivot44 = (main_while_body_bit_concat38_reg < 32'd23);
end
always @(*) begin
		main_NodeBlock41_Pivot42 = (main_while_body_bit_concat38_reg < 32'd35);
end
always @(*) begin
		main_LeafBlock37_SwitchLeaf38 = (main_while_body_bit_concat38_reg == 32'd55);
end
always @(*) begin
		main_LeafBlock35_SwitchLeaf36 = (main_while_body_bit_concat38_reg == 32'd35);
end
always @(*) begin
		main_LeafBlock33_SwitchLeaf34 = (main_while_body_bit_concat38_reg == 32'd23);
end
always @(*) begin
		main_NodeBlock31_Pivot32 = (main_while_body_bit_concat38_reg < 32'd19);
end
always @(*) begin
		main_LeafBlock29_SwitchLeaf30 = (main_while_body_bit_concat38_reg == 32'd19);
end
always @(*) begin
		main_LeafBlock27_SwitchLeaf28 = (main_while_body_bit_concat38_reg == 32'd3);
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_if_else_i_27) & (fsm_stall == 1'd0))) begin
		main_sw_default148_i_results_sroa_28_0249_i = 32'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else62_i_30) & (fsm_stall == 1'd0))) begin
		main_sw_default148_i_results_sroa_28_0249_i = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock18_41) & (fsm_stall == 1'd0)) & (main_LeafBlock18_SwitchLeaf19 == 1'd1))) begin
		main_sw_default148_i_results_sroa_28_0249_i = 32'd65536;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock37_47) & (fsm_stall == 1'd0)) & (main_LeafBlock37_SwitchLeaf38 == 1'd0))) begin
		main_sw_default148_i_results_sroa_28_0249_i = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock35_48) & (fsm_stall == 1'd0)) & (main_LeafBlock35_SwitchLeaf36 == 1'd0))) begin
		main_sw_default148_i_results_sroa_28_0249_i = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock33_49) & (fsm_stall == 1'd0)) & (main_LeafBlock33_SwitchLeaf34 == 1'd0))) begin
		main_sw_default148_i_results_sroa_28_0249_i = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock29_51) & (fsm_stall == 1'd0)) & (main_LeafBlock29_SwitchLeaf30 == 1'd0))) begin
		main_sw_default148_i_results_sroa_28_0249_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_LeafBlock27_52) & (fsm_stall == 1'd0)) & (main_LeafBlock27_SwitchLeaf28 == 1'd0))) */ begin
		main_sw_default148_i_results_sroa_28_0249_i = 32'd0;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_if_else_i_27) & (fsm_stall == 1'd0))) begin
		main_sw_default148_i_results_sroa_28_0249_i_reg <= main_sw_default148_i_results_sroa_28_0249_i;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else62_i_30) & (fsm_stall == 1'd0))) begin
		main_sw_default148_i_results_sroa_28_0249_i_reg <= main_sw_default148_i_results_sroa_28_0249_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock18_41) & (fsm_stall == 1'd0)) & (main_LeafBlock18_SwitchLeaf19 == 1'd1))) begin
		main_sw_default148_i_results_sroa_28_0249_i_reg <= main_sw_default148_i_results_sroa_28_0249_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock37_47) & (fsm_stall == 1'd0)) & (main_LeafBlock37_SwitchLeaf38 == 1'd0))) begin
		main_sw_default148_i_results_sroa_28_0249_i_reg <= main_sw_default148_i_results_sroa_28_0249_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock35_48) & (fsm_stall == 1'd0)) & (main_LeafBlock35_SwitchLeaf36 == 1'd0))) begin
		main_sw_default148_i_results_sroa_28_0249_i_reg <= main_sw_default148_i_results_sroa_28_0249_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock33_49) & (fsm_stall == 1'd0)) & (main_LeafBlock33_SwitchLeaf34 == 1'd0))) begin
		main_sw_default148_i_results_sroa_28_0249_i_reg <= main_sw_default148_i_results_sroa_28_0249_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock29_51) & (fsm_stall == 1'd0)) & (main_LeafBlock29_SwitchLeaf30 == 1'd0))) begin
		main_sw_default148_i_results_sroa_28_0249_i_reg <= main_sw_default148_i_results_sroa_28_0249_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock27_52) & (fsm_stall == 1'd0)) & (main_LeafBlock27_SwitchLeaf28 == 1'd0))) begin
		main_sw_default148_i_results_sroa_28_0249_i_reg <= main_sw_default148_i_results_sroa_28_0249_i;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_if_else_i_27) & (fsm_stall == 1'd0))) begin
		main_sw_default148_i_results_sroa_23_0247_i = 8'd1;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else62_i_30) & (fsm_stall == 1'd0))) begin
		main_sw_default148_i_results_sroa_23_0247_i = 8'd1;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock18_41) & (fsm_stall == 1'd0)) & (main_LeafBlock18_SwitchLeaf19 == 1'd1))) begin
		main_sw_default148_i_results_sroa_23_0247_i = 8'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock37_47) & (fsm_stall == 1'd0)) & (main_LeafBlock37_SwitchLeaf38 == 1'd0))) begin
		main_sw_default148_i_results_sroa_23_0247_i = main_NodeBlock43_results_sroa_23_0_i_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock35_48) & (fsm_stall == 1'd0)) & (main_LeafBlock35_SwitchLeaf36 == 1'd0))) begin
		main_sw_default148_i_results_sroa_23_0247_i = main_NodeBlock43_results_sroa_23_0_i_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock33_49) & (fsm_stall == 1'd0)) & (main_LeafBlock33_SwitchLeaf34 == 1'd0))) begin
		main_sw_default148_i_results_sroa_23_0247_i = main_NodeBlock43_results_sroa_23_0_i_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock29_51) & (fsm_stall == 1'd0)) & (main_LeafBlock29_SwitchLeaf30 == 1'd0))) begin
		main_sw_default148_i_results_sroa_23_0247_i = main_NodeBlock43_results_sroa_23_0_i_reg;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_LeafBlock27_52) & (fsm_stall == 1'd0)) & (main_LeafBlock27_SwitchLeaf28 == 1'd0))) */ begin
		main_sw_default148_i_results_sroa_23_0247_i = main_NodeBlock43_results_sroa_23_0_i_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_if_else_i_27) & (fsm_stall == 1'd0))) begin
		main_sw_default148_i_results_sroa_23_0247_i_reg <= main_sw_default148_i_results_sroa_23_0247_i;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else62_i_30) & (fsm_stall == 1'd0))) begin
		main_sw_default148_i_results_sroa_23_0247_i_reg <= main_sw_default148_i_results_sroa_23_0247_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock18_41) & (fsm_stall == 1'd0)) & (main_LeafBlock18_SwitchLeaf19 == 1'd1))) begin
		main_sw_default148_i_results_sroa_23_0247_i_reg <= main_sw_default148_i_results_sroa_23_0247_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock37_47) & (fsm_stall == 1'd0)) & (main_LeafBlock37_SwitchLeaf38 == 1'd0))) begin
		main_sw_default148_i_results_sroa_23_0247_i_reg <= main_sw_default148_i_results_sroa_23_0247_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock35_48) & (fsm_stall == 1'd0)) & (main_LeafBlock35_SwitchLeaf36 == 1'd0))) begin
		main_sw_default148_i_results_sroa_23_0247_i_reg <= main_sw_default148_i_results_sroa_23_0247_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock33_49) & (fsm_stall == 1'd0)) & (main_LeafBlock33_SwitchLeaf34 == 1'd0))) begin
		main_sw_default148_i_results_sroa_23_0247_i_reg <= main_sw_default148_i_results_sroa_23_0247_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock29_51) & (fsm_stall == 1'd0)) & (main_LeafBlock29_SwitchLeaf30 == 1'd0))) begin
		main_sw_default148_i_results_sroa_23_0247_i_reg <= main_sw_default148_i_results_sroa_23_0247_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock27_52) & (fsm_stall == 1'd0)) & (main_LeafBlock27_SwitchLeaf28 == 1'd0))) begin
		main_sw_default148_i_results_sroa_23_0247_i_reg <= main_sw_default148_i_results_sroa_23_0247_i;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_if_else_i_27) & (fsm_stall == 1'd0))) begin
		main_sw_default148_i_results_sroa_14_0241245_i = main_if_else_i_bit_concat35;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else62_i_30) & (fsm_stall == 1'd0))) begin
		main_sw_default148_i_results_sroa_14_0241245_i = main_if_else62_i_bit_concat31;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock18_41) & (fsm_stall == 1'd0)) & (main_LeafBlock18_SwitchLeaf19 == 1'd1))) begin
		main_sw_default148_i_results_sroa_14_0241245_i = main_NodeBlock24_results_sroa_14_0_i_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock37_47) & (fsm_stall == 1'd0)) & (main_LeafBlock37_SwitchLeaf38 == 1'd0))) begin
		main_sw_default148_i_results_sroa_14_0241245_i = main_NodeBlock43_results_sroa_14_0241_i_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock35_48) & (fsm_stall == 1'd0)) & (main_LeafBlock35_SwitchLeaf36 == 1'd0))) begin
		main_sw_default148_i_results_sroa_14_0241245_i = main_NodeBlock43_results_sroa_14_0241_i_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock33_49) & (fsm_stall == 1'd0)) & (main_LeafBlock33_SwitchLeaf34 == 1'd0))) begin
		main_sw_default148_i_results_sroa_14_0241245_i = main_NodeBlock43_results_sroa_14_0241_i_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock29_51) & (fsm_stall == 1'd0)) & (main_LeafBlock29_SwitchLeaf30 == 1'd0))) begin
		main_sw_default148_i_results_sroa_14_0241245_i = main_NodeBlock43_results_sroa_14_0241_i_reg;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_LeafBlock27_52) & (fsm_stall == 1'd0)) & (main_LeafBlock27_SwitchLeaf28 == 1'd0))) */ begin
		main_sw_default148_i_results_sroa_14_0241245_i = main_NodeBlock43_results_sroa_14_0241_i_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_if_else_i_27) & (fsm_stall == 1'd0))) begin
		main_sw_default148_i_results_sroa_14_0241245_i_reg <= main_sw_default148_i_results_sroa_14_0241245_i;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else62_i_30) & (fsm_stall == 1'd0))) begin
		main_sw_default148_i_results_sroa_14_0241245_i_reg <= main_sw_default148_i_results_sroa_14_0241245_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock18_41) & (fsm_stall == 1'd0)) & (main_LeafBlock18_SwitchLeaf19 == 1'd1))) begin
		main_sw_default148_i_results_sroa_14_0241245_i_reg <= main_sw_default148_i_results_sroa_14_0241245_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock37_47) & (fsm_stall == 1'd0)) & (main_LeafBlock37_SwitchLeaf38 == 1'd0))) begin
		main_sw_default148_i_results_sroa_14_0241245_i_reg <= main_sw_default148_i_results_sroa_14_0241245_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock35_48) & (fsm_stall == 1'd0)) & (main_LeafBlock35_SwitchLeaf36 == 1'd0))) begin
		main_sw_default148_i_results_sroa_14_0241245_i_reg <= main_sw_default148_i_results_sroa_14_0241245_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock33_49) & (fsm_stall == 1'd0)) & (main_LeafBlock33_SwitchLeaf34 == 1'd0))) begin
		main_sw_default148_i_results_sroa_14_0241245_i_reg <= main_sw_default148_i_results_sroa_14_0241245_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock29_51) & (fsm_stall == 1'd0)) & (main_LeafBlock29_SwitchLeaf30 == 1'd0))) begin
		main_sw_default148_i_results_sroa_14_0241245_i_reg <= main_sw_default148_i_results_sroa_14_0241245_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock27_52) & (fsm_stall == 1'd0)) & (main_LeafBlock27_SwitchLeaf28 == 1'd0))) begin
		main_sw_default148_i_results_sroa_14_0241245_i_reg <= main_sw_default148_i_results_sroa_14_0241245_i;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock37_47) & (fsm_stall == 1'd0)) & (main_LeafBlock37_SwitchLeaf38 == 1'd1))) begin
		main_NodeBlock78_results_sroa_28_0248_i = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock35_48) & (fsm_stall == 1'd0)) & (main_LeafBlock35_SwitchLeaf36 == 1'd1))) begin
		main_NodeBlock78_results_sroa_28_0248_i = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock33_49) & (fsm_stall == 1'd0)) & (main_LeafBlock33_SwitchLeaf34 == 1'd1))) begin
		main_NodeBlock78_results_sroa_28_0248_i = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock29_51) & (fsm_stall == 1'd0)) & (main_LeafBlock29_SwitchLeaf30 == 1'd1))) begin
		main_NodeBlock78_results_sroa_28_0248_i = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock27_52) & (fsm_stall == 1'd0)) & (main_LeafBlock27_SwitchLeaf28 == 1'd1))) begin
		main_NodeBlock78_results_sroa_28_0248_i = 32'd0;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_sw_default148_i_53) & (fsm_stall == 1'd0))) */ begin
		main_NodeBlock78_results_sroa_28_0248_i = main_sw_default148_i_results_sroa_28_0249_i_reg;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock37_47) & (fsm_stall == 1'd0)) & (main_LeafBlock37_SwitchLeaf38 == 1'd1))) begin
		main_NodeBlock78_results_sroa_28_0248_i_reg <= main_NodeBlock78_results_sroa_28_0248_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock35_48) & (fsm_stall == 1'd0)) & (main_LeafBlock35_SwitchLeaf36 == 1'd1))) begin
		main_NodeBlock78_results_sroa_28_0248_i_reg <= main_NodeBlock78_results_sroa_28_0248_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock33_49) & (fsm_stall == 1'd0)) & (main_LeafBlock33_SwitchLeaf34 == 1'd1))) begin
		main_NodeBlock78_results_sroa_28_0248_i_reg <= main_NodeBlock78_results_sroa_28_0248_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock29_51) & (fsm_stall == 1'd0)) & (main_LeafBlock29_SwitchLeaf30 == 1'd1))) begin
		main_NodeBlock78_results_sroa_28_0248_i_reg <= main_NodeBlock78_results_sroa_28_0248_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock27_52) & (fsm_stall == 1'd0)) & (main_LeafBlock27_SwitchLeaf28 == 1'd1))) begin
		main_NodeBlock78_results_sroa_28_0248_i_reg <= main_NodeBlock78_results_sroa_28_0248_i;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default148_i_53) & (fsm_stall == 1'd0))) begin
		main_NodeBlock78_results_sroa_28_0248_i_reg <= main_NodeBlock78_results_sroa_28_0248_i;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock37_47) & (fsm_stall == 1'd0)) & (main_LeafBlock37_SwitchLeaf38 == 1'd1))) begin
		main_NodeBlock78_results_sroa_23_0246_i = main_NodeBlock43_results_sroa_23_0_i_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock35_48) & (fsm_stall == 1'd0)) & (main_LeafBlock35_SwitchLeaf36 == 1'd1))) begin
		main_NodeBlock78_results_sroa_23_0246_i = main_NodeBlock43_results_sroa_23_0_i_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock33_49) & (fsm_stall == 1'd0)) & (main_LeafBlock33_SwitchLeaf34 == 1'd1))) begin
		main_NodeBlock78_results_sroa_23_0246_i = main_NodeBlock43_results_sroa_23_0_i_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock29_51) & (fsm_stall == 1'd0)) & (main_LeafBlock29_SwitchLeaf30 == 1'd1))) begin
		main_NodeBlock78_results_sroa_23_0246_i = main_NodeBlock43_results_sroa_23_0_i_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock27_52) & (fsm_stall == 1'd0)) & (main_LeafBlock27_SwitchLeaf28 == 1'd1))) begin
		main_NodeBlock78_results_sroa_23_0246_i = main_NodeBlock43_results_sroa_23_0_i_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_sw_default148_i_53) & (fsm_stall == 1'd0))) */ begin
		main_NodeBlock78_results_sroa_23_0246_i = main_sw_default148_i_results_sroa_23_0247_i_reg;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock37_47) & (fsm_stall == 1'd0)) & (main_LeafBlock37_SwitchLeaf38 == 1'd1))) begin
		main_NodeBlock78_results_sroa_23_0246_i_reg <= main_NodeBlock78_results_sroa_23_0246_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock35_48) & (fsm_stall == 1'd0)) & (main_LeafBlock35_SwitchLeaf36 == 1'd1))) begin
		main_NodeBlock78_results_sroa_23_0246_i_reg <= main_NodeBlock78_results_sroa_23_0246_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock33_49) & (fsm_stall == 1'd0)) & (main_LeafBlock33_SwitchLeaf34 == 1'd1))) begin
		main_NodeBlock78_results_sroa_23_0246_i_reg <= main_NodeBlock78_results_sroa_23_0246_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock29_51) & (fsm_stall == 1'd0)) & (main_LeafBlock29_SwitchLeaf30 == 1'd1))) begin
		main_NodeBlock78_results_sroa_23_0246_i_reg <= main_NodeBlock78_results_sroa_23_0246_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock27_52) & (fsm_stall == 1'd0)) & (main_LeafBlock27_SwitchLeaf28 == 1'd1))) begin
		main_NodeBlock78_results_sroa_23_0246_i_reg <= main_NodeBlock78_results_sroa_23_0246_i;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default148_i_53) & (fsm_stall == 1'd0))) begin
		main_NodeBlock78_results_sroa_23_0246_i_reg <= main_NodeBlock78_results_sroa_23_0246_i;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock37_47) & (fsm_stall == 1'd0)) & (main_LeafBlock37_SwitchLeaf38 == 1'd1))) begin
		main_NodeBlock78_results_sroa_14_0241244_i = main_NodeBlock43_results_sroa_14_0241_i_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock35_48) & (fsm_stall == 1'd0)) & (main_LeafBlock35_SwitchLeaf36 == 1'd1))) begin
		main_NodeBlock78_results_sroa_14_0241244_i = main_NodeBlock43_results_sroa_14_0241_i_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock33_49) & (fsm_stall == 1'd0)) & (main_LeafBlock33_SwitchLeaf34 == 1'd1))) begin
		main_NodeBlock78_results_sroa_14_0241244_i = main_NodeBlock43_results_sroa_14_0241_i_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock29_51) & (fsm_stall == 1'd0)) & (main_LeafBlock29_SwitchLeaf30 == 1'd1))) begin
		main_NodeBlock78_results_sroa_14_0241244_i = main_NodeBlock43_results_sroa_14_0241_i_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock27_52) & (fsm_stall == 1'd0)) & (main_LeafBlock27_SwitchLeaf28 == 1'd1))) begin
		main_NodeBlock78_results_sroa_14_0241244_i = main_NodeBlock43_results_sroa_14_0241_i_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_sw_default148_i_53) & (fsm_stall == 1'd0))) */ begin
		main_NodeBlock78_results_sroa_14_0241244_i = main_sw_default148_i_results_sroa_14_0241245_i_reg;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock37_47) & (fsm_stall == 1'd0)) & (main_LeafBlock37_SwitchLeaf38 == 1'd1))) begin
		main_NodeBlock78_results_sroa_14_0241244_i_reg <= main_NodeBlock78_results_sroa_14_0241244_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock35_48) & (fsm_stall == 1'd0)) & (main_LeafBlock35_SwitchLeaf36 == 1'd1))) begin
		main_NodeBlock78_results_sroa_14_0241244_i_reg <= main_NodeBlock78_results_sroa_14_0241244_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock33_49) & (fsm_stall == 1'd0)) & (main_LeafBlock33_SwitchLeaf34 == 1'd1))) begin
		main_NodeBlock78_results_sroa_14_0241244_i_reg <= main_NodeBlock78_results_sroa_14_0241244_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock29_51) & (fsm_stall == 1'd0)) & (main_LeafBlock29_SwitchLeaf30 == 1'd1))) begin
		main_NodeBlock78_results_sroa_14_0241244_i_reg <= main_NodeBlock78_results_sroa_14_0241244_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock27_52) & (fsm_stall == 1'd0)) & (main_LeafBlock27_SwitchLeaf28 == 1'd1))) begin
		main_NodeBlock78_results_sroa_14_0241244_i_reg <= main_NodeBlock78_results_sroa_14_0241244_i;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default148_i_53) & (fsm_stall == 1'd0))) begin
		main_NodeBlock78_results_sroa_14_0241244_i_reg <= main_NodeBlock78_results_sroa_14_0241244_i;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock37_47) & (fsm_stall == 1'd0)) & (main_LeafBlock37_SwitchLeaf38 == 1'd1))) begin
		main_NodeBlock78_results_sroa_26_0_i = 32'd256;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock35_48) & (fsm_stall == 1'd0)) & (main_LeafBlock35_SwitchLeaf36 == 1'd1))) begin
		main_NodeBlock78_results_sroa_26_0_i = 32'd256;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock33_49) & (fsm_stall == 1'd0)) & (main_LeafBlock33_SwitchLeaf34 == 1'd1))) begin
		main_NodeBlock78_results_sroa_26_0_i = 32'd256;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock29_51) & (fsm_stall == 1'd0)) & (main_LeafBlock29_SwitchLeaf30 == 1'd1))) begin
		main_NodeBlock78_results_sroa_26_0_i = 32'd256;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock27_52) & (fsm_stall == 1'd0)) & (main_LeafBlock27_SwitchLeaf28 == 1'd1))) begin
		main_NodeBlock78_results_sroa_26_0_i = 32'd256;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_sw_default148_i_53) & (fsm_stall == 1'd0))) */ begin
		main_NodeBlock78_results_sroa_26_0_i = 32'd0;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock37_47) & (fsm_stall == 1'd0)) & (main_LeafBlock37_SwitchLeaf38 == 1'd1))) begin
		main_NodeBlock78_results_sroa_26_0_i_reg <= main_NodeBlock78_results_sroa_26_0_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock35_48) & (fsm_stall == 1'd0)) & (main_LeafBlock35_SwitchLeaf36 == 1'd1))) begin
		main_NodeBlock78_results_sroa_26_0_i_reg <= main_NodeBlock78_results_sroa_26_0_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock33_49) & (fsm_stall == 1'd0)) & (main_LeafBlock33_SwitchLeaf34 == 1'd1))) begin
		main_NodeBlock78_results_sroa_26_0_i_reg <= main_NodeBlock78_results_sroa_26_0_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock29_51) & (fsm_stall == 1'd0)) & (main_LeafBlock29_SwitchLeaf30 == 1'd1))) begin
		main_NodeBlock78_results_sroa_26_0_i_reg <= main_NodeBlock78_results_sroa_26_0_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock27_52) & (fsm_stall == 1'd0)) & (main_LeafBlock27_SwitchLeaf28 == 1'd1))) begin
		main_NodeBlock78_results_sroa_26_0_i_reg <= main_NodeBlock78_results_sroa_26_0_i;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default148_i_53) & (fsm_stall == 1'd0))) begin
		main_NodeBlock78_results_sroa_26_0_i_reg <= main_NodeBlock78_results_sroa_26_0_i;
	end
end
always @(*) begin
		main_NodeBlock78_bit_select3 = main_NodeBlock78_results_sroa_28_0248_i_reg[16];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_NodeBlock78_54)) begin
		main_NodeBlock78_bit_select3_reg <= main_NodeBlock78_bit_select3;
	end
end
always @(*) begin
		main_NodeBlock78_bit_select1 = main_NodeBlock78_results_sroa_23_0246_i_reg;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_NodeBlock78_54)) begin
		main_NodeBlock78_bit_select1_reg <= main_NodeBlock78_bit_select1;
	end
end
always @(*) begin
		main_NodeBlock78_Pivot79 = (main_while_body_bit_concat38_reg < 32'd51);
end
always @(*) begin
		main_NodeBlock76_Pivot77 = (main_while_body_bit_concat38_reg < 32'd99);
end
always @(*) begin
		main_NodeBlock74_Pivot75 = (main_while_body_bit_concat38_reg < 32'd103);
end
always @(*) begin
		main_NodeBlock72_Pivot73 = (main_while_body_bit_concat38_reg < 32'd111);
end
always @(*) begin
		main_LeafBlock70_SwitchLeaf71 = (main_while_body_bit_concat38_reg == 32'd111);
end
always @(*) begin
		main_LeafBlock68_SwitchLeaf69 = (main_while_body_bit_concat38_reg == 32'd103);
end
always @(*) begin
		main_LeafBlock66_SwitchLeaf67 = (main_while_body_bit_concat38_reg == 32'd99);
end
always @(*) begin
		main_LeafBlock62_SwitchLeaf63 = (main_while_body_bit_concat38_reg == 32'd55);
end
always @(*) begin
		main_LeafBlock60_SwitchLeaf61 = (main_while_body_bit_concat38_reg == 32'd51);
end
always @(*) begin
		main_NodeBlock58_Pivot59 = (main_while_body_bit_concat38_reg < 32'd23);
end
always @(*) begin
		main_NodeBlock56_Pivot57 = (main_while_body_bit_concat38_reg < 32'd35);
end
always @(*) begin
		main_LeafBlock54_SwitchLeaf55 = (main_while_body_bit_concat38_reg == 32'd35);
end
always @(*) begin
		main_LeafBlock52_SwitchLeaf53 = (main_while_body_bit_concat38_reg == 32'd23);
end
always @(*) begin
		main_NodeBlock50_Pivot51 = (main_while_body_bit_concat38_reg < 32'd19);
end
always @(*) begin
		main_LeafBlock48_SwitchLeaf49 = (main_while_body_bit_concat38_reg == 32'd19);
end
always @(*) begin
		main_LeafBlock46_SwitchLeaf47 = (main_while_body_bit_concat38_reg == 32'd3);
end
always @(*) begin
		main_NodeBlock89_Pivot90 = ($signed($signed({{25{main_while_body_shr6_i_reg[6]}},main_while_body_shr6_i_reg})) < $signed({29'd0,main_NodeBlock89_Pivot90_op1_temp}));
end
always @(*) begin
		main_NodeBlock87_Pivot88 = ($signed($signed({{25{main_while_body_shr6_i_reg[6]}},main_while_body_shr6_i_reg})) < $signed({24'd0,main_NodeBlock87_Pivot88_op1_temp}));
end
always @(*) begin
		main_LeafBlock85_SwitchLeaf86 = ($signed(main_while_body_shr6_i_reg) == 32'd32);
end
always @(*) begin
		main_LeafBlock83_SwitchLeaf84 = ($signed(main_while_body_shr6_i_reg) == 32'd1);
end
always @(*) begin
		main_LeafBlock81_SwitchLeaf82 = ($signed(main_while_body_shr6_i_reg) == 32'd0);
end
always @(*) begin
		main_NodeBlock96_Pivot97 = (main_while_body_bit_concat40_reg < 32'd5);
end
always @(*) begin
		main_LeafBlock94_SwitchLeaf95 = (main_while_body_bit_concat40_reg == 32'd5);
end
always @(*) begin
		main_LeafBlock92_SwitchLeaf93 = (main_while_body_bit_concat40_reg == 32'd0);
end
always @(*) begin
		main_NodeBlock115_Pivot116 = (main_while_body_bit_concat40_reg < 32'd4);
end
always @(*) begin
		main_NodeBlock113_Pivot114 = (main_while_body_bit_concat40_reg < 32'd6);
end
always @(*) begin
		main_NodeBlock111_Pivot112 = (main_while_body_bit_concat40_reg == 32'd7);
end
always @(*) begin
		main_NodeBlock107_Pivot108 = (main_while_body_bit_concat40_reg < 32'd5);
end
always @(*) begin
		main_NodeBlock105_Pivot106 = (main_while_body_bit_concat40_reg < 32'd2);
end
always @(*) begin
		main_NodeBlock103_Pivot104 = (main_while_body_bit_concat40_reg < 32'd3);
end
always @(*) begin
		main_NodeBlock103_1 = (main_NodeBlock103_Pivot104 ? 32'd5 : 32'd6);
end
always @(*) begin
		main_NodeBlock101_Pivot102 = (main_while_body_bit_concat40_reg == 32'd0);
end
always @(*) begin
		main_NodeBlock122_Pivot123 = ($signed($signed({{25{main_while_body_shr6_i_reg[6]}},main_while_body_shr6_i_reg})) < $signed({24'd0,main_NodeBlock122_Pivot123_op1_temp}));
end
always @(*) begin
		main_LeafBlock120_SwitchLeaf121 = ($signed(main_while_body_shr6_i_reg) == 32'd32);
end
always @(*) begin
		main_LeafBlock118_SwitchLeaf119 = ($signed(main_while_body_shr6_i_reg) == 32'd0);
end
always @(*) begin
		main_switch_lookup_i_switch_gep_i = (1'd0 + (4 * main_while_body_bit_concat40_reg));
end
always @(*) begin
		main_switch_lookup_i_switch_load_i = switch_table_out_a;
end
always @(*) begin
		main_switch_lookup54_i_switch_gep56_i = (1'd0 + (4 * main_while_body_bit_concat40_reg));
end
always @(*) begin
		main_switch_lookup54_i_switch_load57_i = switch_table1_out_a;
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock70_58) & (fsm_stall == 1'd0)) & (main_LeafBlock70_SwitchLeaf71 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock68_59) & (fsm_stall == 1'd0)) & (main_LeafBlock68_SwitchLeaf69 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock62_62) & (fsm_stall == 1'd0)) & (main_LeafBlock62_SwitchLeaf63 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock54_66) & (fsm_stall == 1'd0)) & (main_LeafBlock54_SwitchLeaf55 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock52_67) & (fsm_stall == 1'd0)) & (main_LeafBlock52_SwitchLeaf53 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock46_70) & (fsm_stall == 1'd0)) & (main_LeafBlock46_SwitchLeaf47 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock83_74) & (fsm_stall == 1'd0)) & (main_LeafBlock83_SwitchLeaf84 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock94_77) & (fsm_stall == 1'd0)) & (main_LeafBlock94_SwitchLeaf95 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock92_78) & (fsm_stall == 1'd0)) & (main_LeafBlock92_SwitchLeaf93 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default13_i_79) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default16_i_80) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if ((((cur_state == LEGUP_F_main_BB_NodeBlock111_83) & (fsm_stall == 1'd0)) & (main_NodeBlock111_Pivot112 == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock109_84) & (fsm_stall == 1'd0)) & (1'd1 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if ((((cur_state == LEGUP_F_main_BB_NodeBlock107_86) & (fsm_stall == 1'd0)) & (main_NodeBlock107_Pivot108 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if (((cur_state == LEGUP_F_main_BB_NodeBlock103_88) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if ((((cur_state == LEGUP_F_main_BB_NodeBlock101_89) & (fsm_stall == 1'd0)) & (main_NodeBlock101_Pivot102 == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock99_90) & (fsm_stall == 1'd0)) & (1'd1 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock120_93) & (fsm_stall == 1'd0)) & (main_LeafBlock120_SwitchLeaf121 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock118_94) & (fsm_stall == 1'd0)) & (main_LeafBlock118_SwitchLeaf119 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default29_i_95) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default31_i_96) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default48_i_97) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else if (((cur_state == LEGUP_F_main_BB_switch_lookup_i_99) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd256;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_switch_lookup54_i_101) & (fsm_stall == 1'd0))) */ begin
		main_aluDecode_exit_results_sroa_37_0_i6 = 16'd0;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock70_58) & (fsm_stall == 1'd0)) & (main_LeafBlock70_SwitchLeaf71 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock68_59) & (fsm_stall == 1'd0)) & (main_LeafBlock68_SwitchLeaf69 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock62_62) & (fsm_stall == 1'd0)) & (main_LeafBlock62_SwitchLeaf63 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock54_66) & (fsm_stall == 1'd0)) & (main_LeafBlock54_SwitchLeaf55 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock52_67) & (fsm_stall == 1'd0)) & (main_LeafBlock52_SwitchLeaf53 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock46_70) & (fsm_stall == 1'd0)) & (main_LeafBlock46_SwitchLeaf47 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock83_74) & (fsm_stall == 1'd0)) & (main_LeafBlock83_SwitchLeaf84 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock94_77) & (fsm_stall == 1'd0)) & (main_LeafBlock94_SwitchLeaf95 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock92_78) & (fsm_stall == 1'd0)) & (main_LeafBlock92_SwitchLeaf93 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default13_i_79) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default16_i_80) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock111_83) & (fsm_stall == 1'd0)) & (main_NodeBlock111_Pivot112 == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock109_84) & (fsm_stall == 1'd0)) & (1'd1 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock107_86) & (fsm_stall == 1'd0)) & (main_NodeBlock107_Pivot108 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if (((cur_state == LEGUP_F_main_BB_NodeBlock103_88) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock101_89) & (fsm_stall == 1'd0)) & (main_NodeBlock101_Pivot102 == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock99_90) & (fsm_stall == 1'd0)) & (1'd1 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock120_93) & (fsm_stall == 1'd0)) & (main_LeafBlock120_SwitchLeaf121 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock118_94) & (fsm_stall == 1'd0)) & (main_LeafBlock118_SwitchLeaf119 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default29_i_95) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default31_i_96) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default48_i_97) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if (((cur_state == LEGUP_F_main_BB_switch_lookup_i_99) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
	if (((cur_state == LEGUP_F_main_BB_switch_lookup54_i_101) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_37_0_i6_reg <= main_aluDecode_exit_results_sroa_37_0_i6;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock70_58) & (fsm_stall == 1'd0)) & (main_LeafBlock70_SwitchLeaf71 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock68_59) & (fsm_stall == 1'd0)) & (main_LeafBlock68_SwitchLeaf69 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock62_62) & (fsm_stall == 1'd0)) & (main_LeafBlock62_SwitchLeaf63 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock54_66) & (fsm_stall == 1'd0)) & (main_LeafBlock54_SwitchLeaf55 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd16777216;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock52_67) & (fsm_stall == 1'd0)) & (main_LeafBlock52_SwitchLeaf53 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock46_70) & (fsm_stall == 1'd0)) & (main_LeafBlock46_SwitchLeaf47 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock83_74) & (fsm_stall == 1'd0)) & (main_LeafBlock83_SwitchLeaf84 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock94_77) & (fsm_stall == 1'd0)) & (main_LeafBlock94_SwitchLeaf95 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock92_78) & (fsm_stall == 1'd0)) & (main_LeafBlock92_SwitchLeaf93 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default13_i_79) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default16_i_80) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_NodeBlock111_83) & (fsm_stall == 1'd0)) & (main_NodeBlock111_Pivot112 == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock109_84) & (fsm_stall == 1'd0)) & (1'd1 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_NodeBlock107_86) & (fsm_stall == 1'd0)) & (main_NodeBlock107_Pivot108 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_NodeBlock103_88) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_NodeBlock101_89) & (fsm_stall == 1'd0)) & (main_NodeBlock101_Pivot102 == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock99_90) & (fsm_stall == 1'd0)) & (1'd1 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock120_93) & (fsm_stall == 1'd0)) & (main_LeafBlock120_SwitchLeaf121 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock118_94) & (fsm_stall == 1'd0)) & (main_LeafBlock118_SwitchLeaf119 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default29_i_95) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default31_i_96) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default48_i_97) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_switch_lookup_i_99) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_switch_lookup54_i_101) & (fsm_stall == 1'd0))) */ begin
		main_aluDecode_exit_results_sroa_31_0250_i4 = 32'd0;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock70_58) & (fsm_stall == 1'd0)) & (main_LeafBlock70_SwitchLeaf71 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock68_59) & (fsm_stall == 1'd0)) & (main_LeafBlock68_SwitchLeaf69 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock62_62) & (fsm_stall == 1'd0)) & (main_LeafBlock62_SwitchLeaf63 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock54_66) & (fsm_stall == 1'd0)) & (main_LeafBlock54_SwitchLeaf55 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock52_67) & (fsm_stall == 1'd0)) & (main_LeafBlock52_SwitchLeaf53 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock46_70) & (fsm_stall == 1'd0)) & (main_LeafBlock46_SwitchLeaf47 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock83_74) & (fsm_stall == 1'd0)) & (main_LeafBlock83_SwitchLeaf84 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock94_77) & (fsm_stall == 1'd0)) & (main_LeafBlock94_SwitchLeaf95 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock92_78) & (fsm_stall == 1'd0)) & (main_LeafBlock92_SwitchLeaf93 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default13_i_79) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default16_i_80) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock111_83) & (fsm_stall == 1'd0)) & (main_NodeBlock111_Pivot112 == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock109_84) & (fsm_stall == 1'd0)) & (1'd1 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock107_86) & (fsm_stall == 1'd0)) & (main_NodeBlock107_Pivot108 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if (((cur_state == LEGUP_F_main_BB_NodeBlock103_88) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock101_89) & (fsm_stall == 1'd0)) & (main_NodeBlock101_Pivot102 == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock99_90) & (fsm_stall == 1'd0)) & (1'd1 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock120_93) & (fsm_stall == 1'd0)) & (main_LeafBlock120_SwitchLeaf121 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock118_94) & (fsm_stall == 1'd0)) & (main_LeafBlock118_SwitchLeaf119 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default29_i_95) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default31_i_96) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default48_i_97) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if (((cur_state == LEGUP_F_main_BB_switch_lookup_i_99) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
	if (((cur_state == LEGUP_F_main_BB_switch_lookup54_i_101) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_31_0250_i4_reg <= main_aluDecode_exit_results_sroa_31_0250_i4;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock70_58) & (fsm_stall == 1'd0)) & (main_LeafBlock70_SwitchLeaf71 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock68_59) & (fsm_stall == 1'd0)) & (main_LeafBlock68_SwitchLeaf69 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock62_62) & (fsm_stall == 1'd0)) & (main_LeafBlock62_SwitchLeaf63 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock54_66) & (fsm_stall == 1'd0)) & (main_LeafBlock54_SwitchLeaf55 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock52_67) & (fsm_stall == 1'd0)) & (main_LeafBlock52_SwitchLeaf53 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock46_70) & (fsm_stall == 1'd0)) & (main_LeafBlock46_SwitchLeaf47 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd1;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock83_74) & (fsm_stall == 1'd0)) & (main_LeafBlock83_SwitchLeaf84 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock94_77) & (fsm_stall == 1'd0)) & (main_LeafBlock94_SwitchLeaf95 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock92_78) & (fsm_stall == 1'd0)) & (main_LeafBlock92_SwitchLeaf93 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default13_i_79) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default16_i_80) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_NodeBlock111_83) & (fsm_stall == 1'd0)) & (main_NodeBlock111_Pivot112 == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock109_84) & (fsm_stall == 1'd0)) & (1'd1 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_NodeBlock107_86) & (fsm_stall == 1'd0)) & (main_NodeBlock107_Pivot108 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_NodeBlock103_88) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_NodeBlock101_89) & (fsm_stall == 1'd0)) & (main_NodeBlock101_Pivot102 == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock99_90) & (fsm_stall == 1'd0)) & (1'd1 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock120_93) & (fsm_stall == 1'd0)) & (main_LeafBlock120_SwitchLeaf121 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock118_94) & (fsm_stall == 1'd0)) & (main_LeafBlock118_SwitchLeaf119 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default29_i_95) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default31_i_96) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default48_i_97) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_switch_lookup_i_99) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_switch_lookup54_i_101) & (fsm_stall == 1'd0))) */ begin
		main_aluDecode_exit_results_sroa_34_0252_i2 = 16'd0;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock70_58) & (fsm_stall == 1'd0)) & (main_LeafBlock70_SwitchLeaf71 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock68_59) & (fsm_stall == 1'd0)) & (main_LeafBlock68_SwitchLeaf69 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock62_62) & (fsm_stall == 1'd0)) & (main_LeafBlock62_SwitchLeaf63 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock54_66) & (fsm_stall == 1'd0)) & (main_LeafBlock54_SwitchLeaf55 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock52_67) & (fsm_stall == 1'd0)) & (main_LeafBlock52_SwitchLeaf53 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock46_70) & (fsm_stall == 1'd0)) & (main_LeafBlock46_SwitchLeaf47 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock83_74) & (fsm_stall == 1'd0)) & (main_LeafBlock83_SwitchLeaf84 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock94_77) & (fsm_stall == 1'd0)) & (main_LeafBlock94_SwitchLeaf95 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock92_78) & (fsm_stall == 1'd0)) & (main_LeafBlock92_SwitchLeaf93 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default13_i_79) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default16_i_80) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock111_83) & (fsm_stall == 1'd0)) & (main_NodeBlock111_Pivot112 == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock109_84) & (fsm_stall == 1'd0)) & (1'd1 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock107_86) & (fsm_stall == 1'd0)) & (main_NodeBlock107_Pivot108 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if (((cur_state == LEGUP_F_main_BB_NodeBlock103_88) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock101_89) & (fsm_stall == 1'd0)) & (main_NodeBlock101_Pivot102 == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock99_90) & (fsm_stall == 1'd0)) & (1'd1 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock120_93) & (fsm_stall == 1'd0)) & (main_LeafBlock120_SwitchLeaf121 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock118_94) & (fsm_stall == 1'd0)) & (main_LeafBlock118_SwitchLeaf119 == 1'd1))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default29_i_95) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default31_i_96) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default48_i_97) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if (((cur_state == LEGUP_F_main_BB_switch_lookup_i_99) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
	if (((cur_state == LEGUP_F_main_BB_switch_lookup54_i_101) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_results_sroa_34_0252_i2_reg <= main_aluDecode_exit_results_sroa_34_0252_i2;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock70_58) & (fsm_stall == 1'd0)) & (main_LeafBlock70_SwitchLeaf71 == 1'd1))) begin
		main_aluDecode_exit_call13 = 32'd18;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock68_59) & (fsm_stall == 1'd0)) & (main_LeafBlock68_SwitchLeaf69 == 1'd1))) begin
		main_aluDecode_exit_call13 = 32'd19;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock62_62) & (fsm_stall == 1'd0)) & (main_LeafBlock62_SwitchLeaf63 == 1'd1))) begin
		main_aluDecode_exit_call13 = 32'd14;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock54_66) & (fsm_stall == 1'd0)) & (main_LeafBlock54_SwitchLeaf55 == 1'd1))) begin
		main_aluDecode_exit_call13 = 32'd17;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock52_67) & (fsm_stall == 1'd0)) & (main_LeafBlock52_SwitchLeaf53 == 1'd1))) begin
		main_aluDecode_exit_call13 = 32'd15;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock46_70) & (fsm_stall == 1'd0)) & (main_LeafBlock46_SwitchLeaf47 == 1'd1))) begin
		main_aluDecode_exit_call13 = 32'd16;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock83_74) & (fsm_stall == 1'd0)) & (main_LeafBlock83_SwitchLeaf84 == 1'd1))) begin
		main_aluDecode_exit_call13 = 32'd13;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock94_77) & (fsm_stall == 1'd0)) & (main_LeafBlock94_SwitchLeaf95 == 1'd1))) begin
		main_aluDecode_exit_call13 = 32'd7;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock92_78) & (fsm_stall == 1'd0)) & (main_LeafBlock92_SwitchLeaf93 == 1'd1))) begin
		main_aluDecode_exit_call13 = 32'd1;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default13_i_79) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_call13 = 32'd31;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default16_i_80) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_call13 = 32'd31;
	end
	else if ((((cur_state == LEGUP_F_main_BB_NodeBlock111_83) & (fsm_stall == 1'd0)) & (main_NodeBlock111_Pivot112 == 1'd0))) begin
		main_aluDecode_exit_call13 = 32'd3;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock109_84) & (fsm_stall == 1'd0)) & (1'd1 == 1'd1))) begin
		main_aluDecode_exit_call13 = 32'd2;
	end
	else if ((((cur_state == LEGUP_F_main_BB_NodeBlock107_86) & (fsm_stall == 1'd0)) & (main_NodeBlock107_Pivot108 == 1'd1))) begin
		main_aluDecode_exit_call13 = main_while_body_bit_concat40_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_NodeBlock103_88) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_call13 = {29'd0,main_NodeBlock103_1};
	end
	else if ((((cur_state == LEGUP_F_main_BB_NodeBlock101_89) & (fsm_stall == 1'd0)) & (main_NodeBlock101_Pivot102 == 1'd0))) begin
		main_aluDecode_exit_call13 = 32'd12;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock99_90) & (fsm_stall == 1'd0)) & (1'd1 == 1'd1))) begin
		main_aluDecode_exit_call13 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock120_93) & (fsm_stall == 1'd0)) & (main_LeafBlock120_SwitchLeaf121 == 1'd1))) begin
		main_aluDecode_exit_call13 = 32'd8;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock118_94) & (fsm_stall == 1'd0)) & (main_LeafBlock118_SwitchLeaf119 == 1'd1))) begin
		main_aluDecode_exit_call13 = 32'd10;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default29_i_95) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_call13 = 32'd31;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default31_i_96) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_call13 = 0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_default48_i_97) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_call13 = 32'd31;
	end
	else if (((cur_state == LEGUP_F_main_BB_switch_lookup_i_99) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_call13 = main_switch_lookup_i_switch_load_i;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_switch_lookup54_i_101) & (fsm_stall == 1'd0))) */ begin
		main_aluDecode_exit_call13 = main_switch_lookup54_i_switch_load57_i;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock70_58) & (fsm_stall == 1'd0)) & (main_LeafBlock70_SwitchLeaf71 == 1'd1))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock68_59) & (fsm_stall == 1'd0)) & (main_LeafBlock68_SwitchLeaf69 == 1'd1))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock62_62) & (fsm_stall == 1'd0)) & (main_LeafBlock62_SwitchLeaf63 == 1'd1))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock54_66) & (fsm_stall == 1'd0)) & (main_LeafBlock54_SwitchLeaf55 == 1'd1))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock52_67) & (fsm_stall == 1'd0)) & (main_LeafBlock52_SwitchLeaf53 == 1'd1))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock46_70) & (fsm_stall == 1'd0)) & (main_LeafBlock46_SwitchLeaf47 == 1'd1))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock83_74) & (fsm_stall == 1'd0)) & (main_LeafBlock83_SwitchLeaf84 == 1'd1))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock94_77) & (fsm_stall == 1'd0)) & (main_LeafBlock94_SwitchLeaf95 == 1'd1))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock92_78) & (fsm_stall == 1'd0)) & (main_LeafBlock92_SwitchLeaf93 == 1'd1))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default13_i_79) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default16_i_80) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock111_83) & (fsm_stall == 1'd0)) & (main_NodeBlock111_Pivot112 == 1'd0))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock109_84) & (fsm_stall == 1'd0)) & (1'd1 == 1'd1))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock107_86) & (fsm_stall == 1'd0)) & (main_NodeBlock107_Pivot108 == 1'd1))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if (((cur_state == LEGUP_F_main_BB_NodeBlock103_88) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock101_89) & (fsm_stall == 1'd0)) & (main_NodeBlock101_Pivot102 == 1'd0))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock99_90) & (fsm_stall == 1'd0)) & (1'd1 == 1'd1))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock120_93) & (fsm_stall == 1'd0)) & (main_LeafBlock120_SwitchLeaf121 == 1'd1))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock118_94) & (fsm_stall == 1'd0)) & (main_LeafBlock118_SwitchLeaf119 == 1'd1))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default29_i_95) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default31_i_96) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_default48_i_97) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if (((cur_state == LEGUP_F_main_BB_switch_lookup_i_99) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
	if (((cur_state == LEGUP_F_main_BB_switch_lookup54_i_101) & (fsm_stall == 1'd0))) begin
		main_aluDecode_exit_call13_reg <= main_aluDecode_exit_call13;
	end
end
always @(*) begin
		main_aluDecode_exit_arrayidx24 = (1'd0 + (4 * main_while_body_bit_concat45_reg));
end
always @(*) begin
		main_aluDecode_exit_2 = main_while_body_lr_ph_registers_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_aluDecode_exit_103)) begin
		main_aluDecode_exit_2_reg <= main_aluDecode_exit_2;
	end
end
always @(*) begin
		main_aluDecode_exit_tobool = (main_NodeBlock78_results_sroa_26_0_i_reg == 32'd0);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_aluDecode_exit_102)) begin
		main_aluDecode_exit_tobool_reg <= main_aluDecode_exit_tobool;
	end
end
always @(*) begin
		main_if_else_arrayidx27 = (1'd0 + (4 * main_while_body_bit_concat43_reg));
end
always @(*) begin
		main_if_else_3 = main_while_body_lr_ph_registers_out_a;
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_aluDecode_exit_103) & (fsm_stall == 1'd0)) & (main_aluDecode_exit_tobool_reg == 1'd0))) begin
		main_NodeBlock175_aluB_0 = main_NodeBlock78_results_sroa_14_0241244_i_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_if_else_105) & (fsm_stall == 1'd0))) */ begin
		main_NodeBlock175_aluB_0 = main_if_else_3;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_aluDecode_exit_103) & (fsm_stall == 1'd0)) & (main_aluDecode_exit_tobool_reg == 1'd0))) begin
		main_NodeBlock175_aluB_0_reg <= main_NodeBlock175_aluB_0;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else_105) & (fsm_stall == 1'd0))) begin
		main_NodeBlock175_aluB_0_reg <= main_NodeBlock175_aluB_0;
	end
end
always @(*) begin
		main_NodeBlock175_Pivot176 = ($signed(main_aluDecode_exit_call13_reg) < $signed({26'd0,main_NodeBlock175_Pivot176_op1_temp}));
end
always @(*) begin
		main_NodeBlock173_Pivot174 = ($signed(main_aluDecode_exit_call13_reg) < $signed({25'd0,main_NodeBlock173_Pivot174_op1_temp}));
end
always @(*) begin
		main_NodeBlock171_Pivot172 = ($signed(main_aluDecode_exit_call13_reg) < $signed({25'd0,main_NodeBlock171_Pivot172_op1_temp}));
end
always @(*) begin
		main_NodeBlock169_Pivot170 = ($signed(main_aluDecode_exit_call13_reg) < $signed({25'd0,main_NodeBlock169_Pivot170_op1_temp}));
end
always @(*) begin
		main_NodeBlock167_Pivot168 = ($signed(main_aluDecode_exit_call13_reg) < $signed({25'd0,main_NodeBlock167_Pivot168_op1_temp}));
end
always @(*) begin
		main_LeafBlock165_SwitchLeaf166 = (main_aluDecode_exit_call13_reg == 32'd26);
end
always @(*) begin
		main_NodeBlock163_Pivot164 = ($signed(main_aluDecode_exit_call13_reg) < $signed({25'd0,main_NodeBlock163_Pivot164_op1_temp}));
end
always @(*) begin
		main_NodeBlock161_Pivot162 = ($signed(main_aluDecode_exit_call13_reg) < $signed({25'd0,main_NodeBlock161_Pivot162_op1_temp}));
end
always @(*) begin
		main_LeafBlock159_SwitchLeaf160 = (main_aluDecode_exit_call13_reg == 32'd21);
end
always @(*) begin
		main_NodeBlock157_Pivot158 = ($signed(main_aluDecode_exit_call13_reg) < $signed({26'd0,main_NodeBlock157_Pivot158_op1_temp}));
end
always @(*) begin
		main_NodeBlock155_Pivot156 = ($signed(main_aluDecode_exit_call13_reg) < $signed({25'd0,main_NodeBlock155_Pivot156_op1_temp}));
end
always @(*) begin
		main_NodeBlock153_Pivot154 = ($signed(main_aluDecode_exit_call13_reg) < $signed({25'd0,main_NodeBlock153_Pivot154_op1_temp}));
end
always @(*) begin
		main_NodeBlock151_Pivot152 = ($signed(main_aluDecode_exit_call13_reg) < $signed({26'd0,main_NodeBlock151_Pivot152_op1_temp}));
end
always @(*) begin
		main_NodeBlock149_Pivot150 = ($signed(main_aluDecode_exit_call13_reg) < $signed({26'd0,main_NodeBlock149_Pivot150_op1_temp}));
end
always @(*) begin
		main_NodeBlock147_Pivot148 = ($signed(main_aluDecode_exit_call13_reg) < $signed({27'd0,main_NodeBlock147_Pivot148_op1_temp}));
end
always @(*) begin
		main_NodeBlock145_Pivot146 = ($signed(main_aluDecode_exit_call13_reg) < $signed({26'd0,main_NodeBlock145_Pivot146_op1_temp}));
end
always @(*) begin
		main_NodeBlock143_Pivot144 = ($signed(main_aluDecode_exit_call13_reg) < $signed({26'd0,main_NodeBlock143_Pivot144_op1_temp}));
end
always @(*) begin
		main_NodeBlock141_Pivot142 = ($signed(main_aluDecode_exit_call13_reg) < $signed({26'd0,main_NodeBlock141_Pivot142_op1_temp}));
end
always @(*) begin
		main_NodeBlock139_Pivot140 = ($signed(main_aluDecode_exit_call13_reg) < $signed({27'd0,main_NodeBlock139_Pivot140_op1_temp}));
end
always @(*) begin
		main_NodeBlock137_Pivot138 = ($signed(main_aluDecode_exit_call13_reg) < $signed({26'd0,main_NodeBlock137_Pivot138_op1_temp}));
end
always @(*) begin
		main_NodeBlock135_Pivot136 = ($signed(main_aluDecode_exit_call13_reg) < $signed({28'd0,main_NodeBlock135_Pivot136_op1_temp}));
end
always @(*) begin
		main_NodeBlock133_Pivot134 = ($signed(main_aluDecode_exit_call13_reg) < $signed({27'd0,main_NodeBlock133_Pivot134_op1_temp}));
end
always @(*) begin
		main_NodeBlock131_Pivot132 = ($signed(main_aluDecode_exit_call13_reg) < $signed({27'd0,main_NodeBlock131_Pivot132_op1_temp}));
end
always @(*) begin
		main_NodeBlock129_Pivot130 = ($signed(main_aluDecode_exit_call13_reg) < $signed({29'd0,main_NodeBlock129_Pivot130_op1_temp}));
end
always @(*) begin
		main_NodeBlock127_Pivot128 = ($signed(main_aluDecode_exit_call13_reg) < $signed({28'd0,main_NodeBlock127_Pivot128_op1_temp}));
end
always @(*) begin
		main_LeafBlock125_SwitchLeaf126 = (main_aluDecode_exit_call13_reg == 32'd0);
end
always @(*) begin
		main_LeafBlock125_add_i4 = (main_NodeBlock175_aluB_0_reg + main_aluDecode_exit_2_reg);
end
always @(*) begin
		main_LeafBlock125_add_i4_1 = (main_LeafBlock125_SwitchLeaf126 ? main_LeafBlock125_add_i4 : 32'd0);
end
always @(*) begin
		main_sw_bb1_i_sub_i = (main_aluDecode_exit_2_reg - main_NodeBlock175_aluB_0_reg);
end
always @(*) begin
		main_sw_bb5_i_and_i6 = (main_NodeBlock175_aluB_0_reg & main_aluDecode_exit_2_reg);
end
always @(*) begin
		main_sw_bb9_i_or_i = (main_NodeBlock175_aluB_0_reg | main_aluDecode_exit_2_reg);
end
always @(*) begin
		main_sw_bb13_i_xor_i = (main_NodeBlock175_aluB_0_reg ^ main_aluDecode_exit_2_reg);
end
always @(*) begin
		main_sw_bb17_i_cmp_i7 = ($signed(main_aluDecode_exit_2_reg) < $signed(main_NodeBlock175_aluB_0_reg));
end
always @(*) begin
		main_sw_bb17_i_bit_concat12 = {main_sw_bb17_i_bit_concat12_bit_select_operand_0[30:0], main_sw_bb17_i_cmp_i7};
end
always @(*) begin
		main_sw_bb22_i_cmp23_i = (main_aluDecode_exit_2_reg < main_NodeBlock175_aluB_0_reg);
end
always @(*) begin
		main_sw_bb22_i_bit_concat11 = {main_sw_bb22_i_bit_concat11_bit_select_operand_0[30:0], main_sw_bb22_i_cmp23_i};
end
always @(*) begin
		main_sw_bb31_i_shr33_i = ($signed(main_aluDecode_exit_2_reg) >>> main_NodeBlock175_aluB_0_reg);
end
always @(*) begin
		main_sw_bb37_i_shr38_i = ($signed(main_aluDecode_exit_2_reg) >>> main_while_body_bit_concat43_reg);
end
always @(*) begin
		main_sw_bb42_i_shr45_i = (main_aluDecode_exit_2_reg >>> (main_NodeBlock175_aluB_0_reg % 32));
end
always @(*) begin
		main_sw_bb49_i_shr50_i = (main_aluDecode_exit_2_reg >>> (main_while_body_bit_concat43_reg % 32));
end
always @(*) begin
		main_sw_bb54_i_shl_i = (main_aluDecode_exit_2_reg <<< (main_NodeBlock175_aluB_0_reg % 32));
end
always @(*) begin
		main_sw_bb60_i_shl61_i = (main_aluDecode_exit_2_reg <<< (main_while_body_bit_concat43_reg % 32));
end
always @(*) begin
	main_sw_bb65_i_mul_i = main_sw_bb65_i_mul_i_stage0_reg;
end
always @(*) begin
		main_sw_bb73_i_add74_i = (main_NodeBlock175_aluB_0_reg + main_while_body_nextInst_099_reg);
end
always @(*) begin
		main_sw_bb83_i_add84_i = (main_while_body_nextInst_099_reg + 32'd4);
end
always @(*) begin
		main_sw_bb88_i_cmp90_i = (main_aluDecode_exit_2_reg == main_NodeBlock175_aluB_0_reg);
end
always @(*) begin
		main_sw_bb88_i_bit_concat10 = {main_sw_bb88_i_bit_concat10_bit_select_operand_0[6:0], main_sw_bb88_i_cmp90_i};
end
always @(*) begin
		main_sw_bb97_i_not_cmp99_i = (main_aluDecode_exit_2_reg != main_NodeBlock175_aluB_0_reg);
end
always @(*) begin
		main_sw_bb97_i_bit_concat9 = {main_sw_bb97_i_bit_concat9_bit_select_operand_0[6:0], main_sw_bb97_i_not_cmp99_i};
end
always @(*) begin
		main_sw_bb106_i_cmp108_i = ($signed(main_aluDecode_exit_2_reg) < $signed(main_NodeBlock175_aluB_0_reg));
end
always @(*) begin
		main_sw_bb106_i_bit_concat8 = {main_sw_bb106_i_bit_concat8_bit_select_operand_0[6:0], main_sw_bb106_i_cmp108_i};
end
always @(*) begin
		main_sw_bb115_i_not_cmp117_i = ($signed(main_aluDecode_exit_2_reg) >= $signed(main_NodeBlock175_aluB_0_reg));
end
always @(*) begin
		main_sw_bb115_i_bit_concat7 = {main_sw_bb115_i_bit_concat7_bit_select_operand_0[6:0], main_sw_bb115_i_not_cmp117_i};
end
always @(*) begin
		main_sw_bb124_i_cmp126_i = (main_aluDecode_exit_2_reg < main_NodeBlock175_aluB_0_reg);
end
always @(*) begin
		main_sw_bb124_i_bit_concat6 = {main_sw_bb124_i_bit_concat6_bit_select_operand_0[6:0], main_sw_bb124_i_cmp126_i};
end
always @(*) begin
		main_sw_bb133_i_not_cmp135_i = (main_aluDecode_exit_2_reg >= main_NodeBlock175_aluB_0_reg);
end
always @(*) begin
		main_sw_bb133_i_bit_concat5 = {main_sw_bb133_i_bit_concat5_bit_select_operand_0[6:0], main_sw_bb133_i_not_cmp135_i};
end
always @(*) begin
		main_alu_exit_add79_i = (main_NodeBlock175_aluB_0_reg + main_aluDecode_exit_2_reg);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_alu_exit_154)) begin
		main_alu_exit_add79_i_reg <= main_alu_exit_add79_i;
	end
end
always @(*) begin
		main_alu_exit_tobool34 = (main_aluDecode_exit_results_sroa_31_0250_i4_reg == 32'd0);
end
always @(*) begin
		main_if_then38_arrayidx40 = (1'd0 + (4 * main_while_body_bit_concat43_reg));
end
always @(*) begin
		main_if_then38_4 = main_while_body_lr_ph_registers_out_a;
end
always @(*) begin
		main_if_then38_arrayidx41 = (1'd0 + (4 * main_alu_exit_add79_i_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_then38_155)) begin
		main_if_then38_arrayidx41_reg <= main_if_then38_arrayidx41;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock165_111) & (fsm_stall == 1'd0)) & (main_LeafBlock165_SwitchLeaf166 == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock159_114) & (fsm_stall == 1'd0)) & (main_LeafBlock159_SwitchLeaf160 == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_NodeBlock149_119) & (fsm_stall == 1'd0)) & (main_NodeBlock149_Pivot150 == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = main_NodeBlock175_aluB_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_LeafBlock125_131) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = main_LeafBlock125_add_i4_1;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb1_i_132) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = main_sw_bb1_i_sub_i;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb5_i_133) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = main_sw_bb5_i_and_i6;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb9_i_134) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = main_sw_bb9_i_or_i;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb13_i_135) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = main_sw_bb13_i_xor_i;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb17_i_136) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = main_sw_bb17_i_bit_concat12;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb22_i_137) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = main_sw_bb22_i_bit_concat11;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb31_i_138) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = main_sw_bb31_i_shr33_i;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb37_i_139) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = main_sw_bb37_i_shr38_i;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb42_i_140) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = main_sw_bb42_i_shr45_i;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb49_i_141) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = main_sw_bb49_i_shr50_i;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb54_i_142) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = main_sw_bb54_i_shl_i;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb60_i_143) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = main_sw_bb60_i_shl61_i;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb65_i_145) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = main_sw_bb65_i_mul_i;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb73_i_146) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = main_sw_bb73_i_add74_i;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb83_i_147) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = main_sw_bb83_i_add84_i;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb88_i_148) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = 32'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb97_i_149) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = 32'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb106_i_150) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = 32'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb115_i_151) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = 32'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb124_i_152) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = 32'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb133_i_153) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_alu_exit_154) & (fsm_stall == 1'd0)) & (main_alu_exit_tobool34 == 1'd1))) begin
		main_if_end42_results_sroa_0_2_i16 = main_alu_exit_add79_i;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_if_then38_157) & (fsm_stall == 1'd0))) */ begin
		main_if_end42_results_sroa_0_2_i16 = main_alu_exit_add79_i_reg;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock165_111) & (fsm_stall == 1'd0)) & (main_LeafBlock165_SwitchLeaf166 == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock159_114) & (fsm_stall == 1'd0)) & (main_LeafBlock159_SwitchLeaf160 == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock149_119) & (fsm_stall == 1'd0)) & (main_NodeBlock149_Pivot150 == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_LeafBlock125_131) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb1_i_132) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb5_i_133) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb9_i_134) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb13_i_135) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb17_i_136) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb22_i_137) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb31_i_138) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb37_i_139) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb42_i_140) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb49_i_141) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb54_i_142) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb60_i_143) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb65_i_145) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb73_i_146) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb83_i_147) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb88_i_148) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb97_i_149) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb106_i_150) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb115_i_151) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb124_i_152) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb133_i_153) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if ((((cur_state == LEGUP_F_main_BB_alu_exit_154) & (fsm_stall == 1'd0)) & (main_alu_exit_tobool34 == 1'd1))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
	if (((cur_state == LEGUP_F_main_BB_if_then38_157) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_0_2_i16_reg <= main_if_end42_results_sroa_0_2_i16;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock165_111) & (fsm_stall == 1'd0)) & (main_LeafBlock165_SwitchLeaf166 == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock159_114) & (fsm_stall == 1'd0)) & (main_LeafBlock159_SwitchLeaf160 == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_NodeBlock149_119) & (fsm_stall == 1'd0)) & (main_NodeBlock149_Pivot150 == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_LeafBlock125_131) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb1_i_132) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb5_i_133) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb9_i_134) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb13_i_135) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb17_i_136) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb22_i_137) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb31_i_138) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb37_i_139) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb42_i_140) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb49_i_141) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb54_i_142) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb60_i_143) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb65_i_145) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb73_i_146) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb83_i_147) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd1;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb88_i_148) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = main_sw_bb88_i_bit_concat10;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb97_i_149) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = main_sw_bb97_i_bit_concat9;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb106_i_150) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = main_sw_bb106_i_bit_concat8;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb115_i_151) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = main_sw_bb115_i_bit_concat7;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb124_i_152) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = main_sw_bb124_i_bit_concat6;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb133_i_153) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15 = main_sw_bb133_i_bit_concat5;
	end
	else if ((((cur_state == LEGUP_F_main_BB_alu_exit_154) & (fsm_stall == 1'd0)) & (main_alu_exit_tobool34 == 1'd1))) begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_if_then38_157) & (fsm_stall == 1'd0))) */ begin
		main_if_end42_results_sroa_53_6_i15 = 8'd0;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock165_111) & (fsm_stall == 1'd0)) & (main_LeafBlock165_SwitchLeaf166 == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock159_114) & (fsm_stall == 1'd0)) & (main_LeafBlock159_SwitchLeaf160 == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock149_119) & (fsm_stall == 1'd0)) & (main_NodeBlock149_Pivot150 == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_LeafBlock125_131) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb1_i_132) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb5_i_133) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb9_i_134) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb13_i_135) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb17_i_136) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb22_i_137) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb31_i_138) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb37_i_139) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb42_i_140) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb49_i_141) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb54_i_142) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb60_i_143) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb65_i_145) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb73_i_146) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb83_i_147) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb88_i_148) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb97_i_149) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb106_i_150) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb115_i_151) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb124_i_152) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb133_i_153) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if ((((cur_state == LEGUP_F_main_BB_alu_exit_154) & (fsm_stall == 1'd0)) & (main_alu_exit_tobool34 == 1'd1))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
	if (((cur_state == LEGUP_F_main_BB_if_then38_157) & (fsm_stall == 1'd0))) begin
		main_if_end42_results_sroa_53_6_i15_reg <= main_if_end42_results_sroa_53_6_i15;
	end
end
always @(*) begin
		main_if_end42_tobool43 = (main_aluDecode_exit_results_sroa_34_0252_i2_reg == 16'd0);
end
always @(*) begin
		main_if_then47_arrayidx49 = (1'd0 + (4 * main_if_end42_results_sroa_0_2_i16_reg));
end
always @(*) begin
		main_if_then47_5 = main_while_body_lr_ph_memory_out_a;
end
always @(*) begin
		main_if_then47_arrayidx50 = (1'd0 + (4 * main_while_body_bit_concat41_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_then47_159)) begin
		main_if_then47_arrayidx50_reg <= main_if_then47_arrayidx50;
	end
end
always @(*) begin
		main_if_else51_tobool52 = (main_aluDecode_exit_results_sroa_37_0_i6_reg == 16'd0);
end
always @(*) begin
		main_if_then56_arrayidx59 = (1'd0 + (4 * main_while_body_bit_concat41_reg));
end
always @(*) begin
		main_if_end61_tobool63 = (main_if_end42_results_sroa_53_6_i15_reg == 8'd0);
end
always @(*) begin
		main_if_end61_bit_concat4 = {{main_if_end61_bit_concat4_bit_select_operand_0[14:0], main_NodeBlock78_bit_select3_reg}, main_if_end61_bit_concat4_bit_select_operand_4[15:0]};
end
always @(*) begin
		main_if_end61_tobool66 = (main_if_end61_bit_concat4 == 32'd0);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end61_165)) begin
		main_if_end61_tobool66_reg <= main_if_end61_tobool66;
	end
end
always @(*) begin
		main_if_then_i1_bit_concat2 = {main_if_then_i1_bit_concat2_bit_select_operand_0[6:0], main_NodeBlock78_bit_select1_reg};
end
always @(*) begin
		main_if_then_i1_tobool65 = (main_if_then_i1_bit_concat2 == 8'd0);
end
always @(*) begin
		main_if_then8_i_add_i = (main_NodeBlock78_results_sroa_14_0241244_i_reg + main_while_body_nextInst_099_reg);
end
always @(*) begin
		main_if_then13_i_add14_i = (main_aluDecode_exit_2_reg + main_NodeBlock78_results_sroa_14_0241244_i_reg);
end
always @(*) begin
		main_if_then13_i_bit_select = main_if_then13_i_add14_i[31:1];
end
always @(*) begin
		main_if_then13_i_bit_concat = {main_if_then13_i_bit_select[30:0], main_if_then13_i_bit_concat_bit_select_operand_2};
end
always @(*) begin
		main_if_else15_i_add16_i = (main_while_body_nextInst_099_reg + 32'd4);
end
always @(*) begin
		main_if_else18_i_add19_i = (main_while_body_nextInst_099_reg + 32'd4);
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_if_then8_i_167) & (fsm_stall == 1'd0))) begin
		main_addressCalculator_exit_newPc_0_i = main_if_then8_i_add_i;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_then13_i_169) & (fsm_stall == 1'd0))) begin
		main_addressCalculator_exit_newPc_0_i = main_if_then13_i_bit_concat;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else15_i_170) & (fsm_stall == 1'd0))) begin
		main_addressCalculator_exit_newPc_0_i = main_if_else15_i_add16_i;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_if_else18_i_171) & (fsm_stall == 1'd0))) */ begin
		main_addressCalculator_exit_newPc_0_i = main_if_else18_i_add19_i;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_if_then8_i_167) & (fsm_stall == 1'd0))) begin
		main_addressCalculator_exit_newPc_0_i_reg <= main_addressCalculator_exit_newPc_0_i;
	end
	if (((cur_state == LEGUP_F_main_BB_if_then13_i_169) & (fsm_stall == 1'd0))) begin
		main_addressCalculator_exit_newPc_0_i_reg <= main_addressCalculator_exit_newPc_0_i;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else15_i_170) & (fsm_stall == 1'd0))) begin
		main_addressCalculator_exit_newPc_0_i_reg <= main_addressCalculator_exit_newPc_0_i;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else18_i_171) & (fsm_stall == 1'd0))) begin
		main_addressCalculator_exit_newPc_0_i_reg <= main_addressCalculator_exit_newPc_0_i;
	end
end
always @(*) begin
		main_addressCalculator_exit_cmp = (main_while_body_1_reg != 32'd0);
end
always @(*) begin
		main_addressCalculator_exit_cmp21 = ($signed(main_while_body_nextInst_099_reg) < $signed({19'd0,main_addressCalculator_exit_cmp21_op1_temp}));
end
always @(*) begin
		main_addressCalculator_exit_or_cond = (main_addressCalculator_exit_cmp & main_addressCalculator_exit_cmp21);
end
always @(*) begin
		main_if_end61_while_body_crit_edge_arrayidx23_phi_ = (1'd0 + (4 * main_addressCalculator_exit_newPc_0_i_reg));
end
always @(*) begin
		main_if_end61_while_body_crit_edge_pre100 = main_while_body_lr_ph_instMemory_out_a;
end
assign main_while_end_arrayidx68_phi_trans_insert = (1'd0 + (4 * 32'd22));
always @(*) begin
		main_while_end_pre = main_while_body_lr_ph_registers_out_a;
end
always @(*) begin
	switch_table_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_switch_lookup_i_98)) begin
		switch_table_address_a = (main_switch_lookup_i_switch_gep_i >>> 3'd2);
	end
end
assign switch_table_address_b = 'dx;
always @(*) begin
	switch_table1_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_switch_lookup54_i_100)) begin
		switch_table1_address_a = (main_switch_lookup54_i_switch_gep56_i >>> 3'd2);
	end
end
assign switch_table1_address_b = 'dx;
always @(*) begin
	main_while_body_lr_ph_registers_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_while_body_i_2)) begin
		main_while_body_lr_ph_registers_address_a = (main_while_body_i_s_010_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_lr_ph_registers_address_a = (main_legup_memset_4_exit_arrayidx22_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_aluDecode_exit_102)) begin
		main_while_body_lr_ph_registers_address_a = (main_aluDecode_exit_arrayidx24 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_else_104)) begin
		main_while_body_lr_ph_registers_address_a = (main_if_else_arrayidx27 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then38_155)) begin
		main_while_body_lr_ph_registers_address_a = (main_if_then38_arrayidx40 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then47_160)) begin
		main_while_body_lr_ph_registers_address_a = (main_if_then47_arrayidx50_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then56_163)) begin
		main_while_body_lr_ph_registers_address_a = (main_if_then56_arrayidx59 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_while_end_175)) begin
		main_while_body_lr_ph_registers_address_a = (main_while_end_arrayidx68_phi_trans_insert >>> 3'd2);
	end
end
always @(*) begin
	main_while_body_lr_ph_registers_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_while_body_i_2)) begin
		main_while_body_lr_ph_registers_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_lr_ph_registers_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then47_160)) begin
		main_while_body_lr_ph_registers_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then56_163)) begin
		main_while_body_lr_ph_registers_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_while_body_lr_ph_registers_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_while_body_i_2)) begin
		main_while_body_lr_ph_registers_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_while_body_15)) begin
		main_while_body_lr_ph_registers_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then47_160)) begin
		main_while_body_lr_ph_registers_in_a = main_if_then47_5;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then56_163)) begin
		main_while_body_lr_ph_registers_in_a = main_if_end42_results_sroa_0_2_i16_reg;
	end
end
always @(*) begin
	main_while_body_lr_ph_instMemory_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_while_body_lr_ph_instMemory_address_a = (main_legup_memset_4_exit_arrayidx >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_5)) begin
		main_while_body_lr_ph_instMemory_address_a = (main_legup_memset_4_exit_arrayidx2_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_6)) begin
		main_while_body_lr_ph_instMemory_address_a = (main_legup_memset_4_exit_arrayidx4_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_7)) begin
		main_while_body_lr_ph_instMemory_address_a = (main_legup_memset_4_exit_arrayidx6_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_8)) begin
		main_while_body_lr_ph_instMemory_address_a = (main_legup_memset_4_exit_arrayidx8_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_9)) begin
		main_while_body_lr_ph_instMemory_address_a = (main_legup_memset_4_exit_arrayidx10_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_10)) begin
		main_while_body_lr_ph_instMemory_address_a = (main_legup_memset_4_exit_arrayidx12_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_11)) begin
		main_while_body_lr_ph_instMemory_address_a = (main_legup_memset_4_exit_arrayidx14_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_12)) begin
		main_while_body_lr_ph_instMemory_address_a = (main_legup_memset_4_exit_arrayidx16_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_13)) begin
		main_while_body_lr_ph_instMemory_address_a = (main_legup_memset_4_exit_arrayidx18_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_end61_while_body_crit_edge_173)) begin
		main_while_body_lr_ph_instMemory_address_a = (main_if_end61_while_body_crit_edge_arrayidx23_phi_ >>> 3'd2);
	end
end
always @(*) begin
	main_while_body_lr_ph_instMemory_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_while_body_lr_ph_instMemory_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_5)) begin
		main_while_body_lr_ph_instMemory_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_6)) begin
		main_while_body_lr_ph_instMemory_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_7)) begin
		main_while_body_lr_ph_instMemory_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_8)) begin
		main_while_body_lr_ph_instMemory_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_9)) begin
		main_while_body_lr_ph_instMemory_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_10)) begin
		main_while_body_lr_ph_instMemory_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_11)) begin
		main_while_body_lr_ph_instMemory_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_12)) begin
		main_while_body_lr_ph_instMemory_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_13)) begin
		main_while_body_lr_ph_instMemory_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_while_body_lr_ph_instMemory_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_while_body_lr_ph_instMemory_in_a = 32'd536871187;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_5)) begin
		main_while_body_lr_ph_instMemory_in_a = 32'd8388847;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_6)) begin
		main_while_body_lr_ph_instMemory_in_a = -32'd8322797;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_7)) begin
		main_while_body_lr_ph_instMemory_in_a = 32'd10559523;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_8)) begin
		main_while_body_lr_ph_instMemory_in_a = 32'd5592163;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_9)) begin
		main_while_body_lr_ph_instMemory_in_a = -32'd719597;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_10)) begin
		main_while_body_lr_ph_instMemory_in_a = 32'd75139;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_11)) begin
		main_while_body_lr_ph_instMemory_in_a = 32'd8388719;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_12)) begin
		main_while_body_lr_ph_instMemory_in_a = 32'd4268163;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_13)) begin
		main_while_body_lr_ph_instMemory_in_a = 32'd32871;
	end
end
always @(*) begin
	main_while_body_lr_ph_instMemory_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_while_body_lr_ph_instMemory_address_b = (main_legup_memset_4_exit_arrayidx1 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_5)) begin
		main_while_body_lr_ph_instMemory_address_b = (main_legup_memset_4_exit_arrayidx3_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_6)) begin
		main_while_body_lr_ph_instMemory_address_b = (main_legup_memset_4_exit_arrayidx5_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_7)) begin
		main_while_body_lr_ph_instMemory_address_b = (main_legup_memset_4_exit_arrayidx7_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_8)) begin
		main_while_body_lr_ph_instMemory_address_b = (main_legup_memset_4_exit_arrayidx9_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_9)) begin
		main_while_body_lr_ph_instMemory_address_b = (main_legup_memset_4_exit_arrayidx11_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_10)) begin
		main_while_body_lr_ph_instMemory_address_b = (main_legup_memset_4_exit_arrayidx13_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_11)) begin
		main_while_body_lr_ph_instMemory_address_b = (main_legup_memset_4_exit_arrayidx15_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_12)) begin
		main_while_body_lr_ph_instMemory_address_b = (main_legup_memset_4_exit_arrayidx17_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_13)) begin
		main_while_body_lr_ph_instMemory_address_b = (main_legup_memset_4_exit_arrayidx19_reg >>> 3'd2);
	end
end
always @(*) begin
	main_while_body_lr_ph_instMemory_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_while_body_lr_ph_instMemory_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_5)) begin
		main_while_body_lr_ph_instMemory_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_6)) begin
		main_while_body_lr_ph_instMemory_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_7)) begin
		main_while_body_lr_ph_instMemory_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_8)) begin
		main_while_body_lr_ph_instMemory_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_9)) begin
		main_while_body_lr_ph_instMemory_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_10)) begin
		main_while_body_lr_ph_instMemory_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_11)) begin
		main_while_body_lr_ph_instMemory_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_12)) begin
		main_while_body_lr_ph_instMemory_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_13)) begin
		main_while_body_lr_ph_instMemory_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_while_body_lr_ph_instMemory_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_4)) begin
		main_while_body_lr_ph_instMemory_in_b = 32'd4195603;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_5)) begin
		main_while_body_lr_ph_instMemory_in_b = 32'd67108975;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_6)) begin
		main_while_body_lr_ph_instMemory_in_b = 32'd1122851;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_7)) begin
		main_while_body_lr_ph_instMemory_in_b = 32'd1049235;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_8)) begin
		main_while_body_lr_ph_instMemory_in_b = 32'd25165935;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_9)) begin
		main_while_body_lr_ph_instMemory_in_b = -32'd27266833;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_10)) begin
		main_while_body_lr_ph_instMemory_in_b = 32'd45417779;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_11)) begin
		main_while_body_lr_ph_instMemory_in_b = 32'd1049875;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_12)) begin
		main_while_body_lr_ph_instMemory_in_b = 32'd8454419;
	end
	if ((cur_state == LEGUP_F_main_BB_legup_memset_4_exit_13)) begin
		main_while_body_lr_ph_instMemory_in_b = 32'd10488627;
	end
end
always @(*) begin
	main_while_body_lr_ph_memory_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_if_then38_156)) begin
		main_while_body_lr_ph_memory_address_a = (main_if_then38_arrayidx41_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then47_159)) begin
		main_while_body_lr_ph_memory_address_a = (main_if_then47_arrayidx49 >>> 3'd2);
	end
end
always @(*) begin
	main_while_body_lr_ph_memory_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_if_then38_156)) begin
		main_while_body_lr_ph_memory_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_while_body_lr_ph_memory_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_if_then38_156)) begin
		main_while_body_lr_ph_memory_in_a = main_if_then38_4;
	end
end
assign main_while_body_bit_concat45_bit_select_operand_0 = 27'd0;
assign main_while_body_bit_concat43_bit_select_operand_0 = 27'd0;
assign main_while_body_bit_concat41_bit_select_operand_0 = 27'd0;
assign main_while_body_bit_concat40_bit_select_operand_0 = 29'd0;
assign main_while_body_bit_concat38_bit_select_operand_0 = 25'd0;
assign main_if_then_i_bit_concat36_bit_select_operand_0 = -21'd2;
assign main_if_then_i_bit_concat36_bit_select_operand_6 = 1'd0;
assign main_if_else_i_bit_concat35_bit_select_operand_2 = 18'd0;
assign main_if_else_i_bit_concat35_bit_select_operand_6 = 1'd0;
assign main_if_else_i_bit_concat35_bit_select_operand_12 = 1'd0;
assign main_if_then44_i_bit_concat33_bit_select_operand_0 = -12'd1;
assign main_if_then44_i_bit_concat33_bit_select_operand_8 = 1'd0;
assign main_if_else62_i_bit_concat31_bit_select_operand_2 = 11'd0;
assign main_if_else62_i_bit_concat31_bit_select_operand_12 = 1'd0;
assign main_if_then88_i_bit_concat26_bit_select_operand_0 = -21'd1;
assign main_if_then88_i_bit_concat26_bit_select_operand_4 = 1'd0;
assign main_sw_epilog_thread242_i_bit_concat22_bit_select_operand_2 = 19'd0;
assign main_sw_epilog_thread242_i_bit_concat22_bit_select_operand_6 = 1'd0;
assign main_sw_bb118_i_bit_concat18_bit_select_operand_2 = 12'd0;
assign main_if_then126_i_bit_concat15_bit_select_operand_0 = -21'd1;
assign main_if_else131_i_bit_concat14_bit_select_operand_0 = 21'd0;
assign main_NodeBlock89_Pivot90_op1_temp = 32'd1;
assign main_NodeBlock87_Pivot88_op1_temp = 32'd32;
assign main_NodeBlock122_Pivot123_op1_temp = 32'd32;
assign main_NodeBlock175_Pivot176_op1_temp = 32'd12;
assign main_NodeBlock173_Pivot174_op1_temp = 32'd20;
assign main_NodeBlock171_Pivot172_op1_temp = 32'd24;
assign main_NodeBlock169_Pivot170_op1_temp = 32'd25;
assign main_NodeBlock167_Pivot168_op1_temp = 32'd26;
assign main_NodeBlock163_Pivot164_op1_temp = 32'd21;
assign main_NodeBlock161_Pivot162_op1_temp = 32'd23;
assign main_NodeBlock157_Pivot158_op1_temp = 32'd15;
assign main_NodeBlock155_Pivot156_op1_temp = 32'd16;
assign main_NodeBlock153_Pivot154_op1_temp = 32'd18;
assign main_NodeBlock151_Pivot152_op1_temp = 32'd13;
assign main_NodeBlock149_Pivot150_op1_temp = 32'd14;
assign main_NodeBlock147_Pivot148_op1_temp = 32'd6;
assign main_NodeBlock145_Pivot146_op1_temp = 32'd9;
assign main_NodeBlock143_Pivot144_op1_temp = 32'd10;
assign main_NodeBlock141_Pivot142_op1_temp = 32'd11;
assign main_NodeBlock139_Pivot140_op1_temp = 32'd7;
assign main_NodeBlock137_Pivot138_op1_temp = 32'd8;
assign main_NodeBlock135_Pivot136_op1_temp = 32'd3;
assign main_NodeBlock133_Pivot134_op1_temp = 32'd4;
assign main_NodeBlock131_Pivot132_op1_temp = 32'd5;
assign main_NodeBlock129_Pivot130_op1_temp = 32'd1;
assign main_NodeBlock127_Pivot128_op1_temp = 32'd2;
assign main_sw_bb17_i_bit_concat12_bit_select_operand_0 = 31'd0;
assign main_sw_bb22_i_bit_concat11_bit_select_operand_0 = 31'd0;
always @(*) begin
	legup_mult_main_sw_bb65_i_mul_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_sw_bb65_i_mul_i_en == 1'd1)) begin
		main_sw_bb65_i_mul_i_stage0_reg <= (main_NodeBlock175_aluB_0_reg * main_aluDecode_exit_2_reg);
	end
end
assign main_sw_bb88_i_bit_concat10_bit_select_operand_0 = 7'd0;
assign main_sw_bb97_i_bit_concat9_bit_select_operand_0 = 7'd0;
assign main_sw_bb106_i_bit_concat8_bit_select_operand_0 = 7'd0;
assign main_sw_bb115_i_bit_concat7_bit_select_operand_0 = 7'd0;
assign main_sw_bb124_i_bit_concat6_bit_select_operand_0 = 7'd0;
assign main_sw_bb133_i_bit_concat5_bit_select_operand_0 = 7'd0;
assign main_if_end61_bit_concat4_bit_select_operand_0 = 15'd0;
assign main_if_end61_bit_concat4_bit_select_operand_4 = 16'd0;
assign main_if_then_i1_bit_concat2_bit_select_operand_0 = 7'd0;
assign main_if_then13_i_bit_concat_bit_select_operand_2 = 1'd0;
assign main_addressCalculator_exit_cmp21_op1_temp = 32'd1024;
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		finish <= 1'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_while_end_176)) begin
		finish <= (fsm_stall == 1'd0);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		return_val <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_while_end_176)) begin
		return_val <= 32'd0;
	end
end

endmodule
module ram_dual_port
(
	clk,
	clken,
	address_a,
	address_b,
	wren_a,
	data_a,
	byteena_a,
	wren_b,
	data_b,
	byteena_b,
	q_b,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  width_b = 1'd0;
parameter  widthad_b = 1'd0;
parameter  numwords_b = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
parameter  width_be_b = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input [(widthad_b-1):0] address_b;
output wire [(width_b-1):0] q_b;
wire [(width_b-1):0] q_b_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
input  wren_b;
input [(width_b-1):0] data_b;
input [width_be_b-1:0] byteena_b;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
	.address_b (address_b),
    .addressstall_b (1'd0),
    .rden_b (clken),
    .q_b (q_b),
    .wren_a (wren_a),
    .data_a (data_a),
    .wren_b (wren_b),
    .data_b (data_b),
    .byteena_b (byteena_b),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.width_byteena_b = width_be_b,
    altsyncram_component.operation_mode = "BIDIR_DUAL_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "CycloneIV",
    altsyncram_component.clock_enable_input_b = "BYPASS",
    altsyncram_component.clock_enable_output_b = "BYPASS",
    altsyncram_component.outdata_aclr_b = "NONE",
    altsyncram_component.outdata_reg_b = output_registered,
    altsyncram_component.numwords_b = numwords_b,
    altsyncram_component.widthad_b = widthad_b,
    altsyncram_component.width_b = width_b,
    altsyncram_component.address_reg_b = "CLOCK0",
    altsyncram_component.byteena_reg_b = "CLOCK0",
    altsyncram_component.indata_reg_b = "CLOCK0",
    altsyncram_component.wrcontrol_wraddress_reg_b = "CLOCK0",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
module ram_single_port_intel
(
	clk,
	clken,
	address_a,
	wren_a,
	data_a,
	byteena_a,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
    .wren_a (wren_a),
    .data_a (data_a),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.operation_mode = "SINGLE_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "CycloneIV",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
module rom_dual_port
(
	clk,
	clken,
	address_a,
	q_a,
	address_b,
	q_b
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  width_b = 1'd0;
parameter  widthad_b = 1'd0;
parameter  numwords_b = 1'd0;
parameter  init_file = {`MEM_INIT_DIR, "UNUSED.mif"};
parameter  latency = 1;

input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
reg [(width_a-1):0] q_a_wire;
input [(widthad_b-1):0] address_b;
output wire [(width_b-1):0] q_b;
reg [(width_b-1):0] q_b_wire;

(* ram_init_file = init_file *) reg [width_a-1:0] ram [numwords_a-1:0];

integer i;
/* synthesis translate_off */
ALTERA_MF_MEMORY_INITIALIZATION mem ();
reg [8*256:1] ram_ver_file;
initial begin
	if (init_file == {`MEM_INIT_DIR, "UNUSED.mif"})
    begin
		for (i = 0; i < numwords_a; i = i + 1)
			ram[i] = 0;
    end
	else
    begin
        // modelsim can't read .mif files directly. So use Altera function to
        // convert them to .ver files
        mem.convert_to_ver_file(init_file, width_a, ram_ver_file);
        $readmemh(ram_ver_file, ram);
    end
end
/* synthesis translate_on */

localparam input_latency = ((latency - 1) >> 1);
localparam output_latency = (latency - 1) - input_latency;
integer j;

reg [(widthad_a-1):0] address_a_reg[input_latency:0];
reg [(widthad_b-1):0] address_b_reg[input_latency:0];

always @(*)
begin
  address_a_reg[0] = address_a;
  address_b_reg[0] = address_b;
end

always @(posedge clk)
if (clken)
begin
   for (j = 0; j < input_latency; j=j+1)
   begin
       address_a_reg[j+1] <= address_a_reg[j];
       address_b_reg[j+1] <= address_b_reg[j];
   end
end

always @ (posedge clk)
if (clken)
begin
    q_a_wire <= ram[address_a_reg[input_latency]];
end

always @ (posedge clk)
if (clken)
begin
    q_b_wire <= ram[address_b_reg[input_latency]];
end


reg [(width_a-1):0] q_a_reg[output_latency:0];

always @(*)
begin
   q_a_reg[0] <= q_a_wire;
end

always @(posedge clk)
if (clken)
begin
   for (j = 0; j < output_latency; j=j+1)
   begin
       q_a_reg[j+1] <= q_a_reg[j];
   end
end

assign q_a = q_a_reg[output_latency];
reg [(width_b-1):0] q_b_reg[output_latency:0];

always @(*)
begin
   q_b_reg[0] <= q_b_wire;
end

always @(posedge clk)
if (clken)
begin
   for (j = 0; j < output_latency; j=j+1)
   begin
       q_b_reg[j+1] <= q_b_reg[j];
   end
end

assign q_b = q_b_reg[output_latency];

endmodule
`timescale 1 ns / 1 ns
module main_tb
(
);

reg  clk;
reg  reset;
reg  start;
wire [31:0] return_val;
wire  finish;


top top_inst (
	.clk (clk),
	.reset (reset),
	.start (start),
	.finish (finish),
	.return_val (return_val)
);




initial 
    clk = 0;
always @(clk)
    clk <= #10 ~clk;

initial begin
//$monitor("At t=%t clk=%b %b %b %b %d", $time, clk, reset, start, finish, return_val);
reset <= 1;
@(negedge clk);
reset <= 0;
start <= 1;
@(negedge clk);
start <= 0;
end

always@(posedge clk) begin
    if (finish == 1) begin
        $display("At t=%t clk=%b finish=%b return_val=%d", $time, clk, finish, return_val);
        $display("Cycles: %d", ($time-50)/20);
        $finish;
    end
end


endmodule
